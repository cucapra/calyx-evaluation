/* verilator lint_off WIDTH */
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule

module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule

module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

// Component Signature
module mac_pe (
      input wire [31:0] top,
      input wire [31:0] left,
      input wire go,
      input wire clk,
      output wire [31:0] down,
      output wire [31:0] right,
      output wire [31:0] out,
      output wire done
  );
  
  // Structure wire declarations
  wire [31:0] mul_left;
  wire [31:0] mul_right;
  wire mul_go;
  wire mul_clk;
  wire [31:0] mul_out;
  wire mul_done;
  wire [31:0] add_left;
  wire [31:0] add_right;
  wire [31:0] add_out;
  wire [31:0] mul_reg_in;
  wire mul_reg_write_en;
  wire mul_reg_clk;
  wire [31:0] mul_reg_out;
  wire mul_reg_done;
  wire [31:0] acc_in;
  wire acc_write_en;
  wire acc_clk;
  wire [31:0] acc_out;
  wire acc_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_mult_pipe #(32) mul (
      .left(mul_left),
      .right(mul_right),
      .go(mul_go),
      .clk(clk),
      .out(mul_out),
      .done(mul_done)
  );
  
  std_add #(32) add (
      .left(add_left),
      .right(add_right),
      .out(add_out)
  );
  
  std_reg #(32) mul_reg (
      .in(mul_reg_in),
      .write_en(mul_reg_write_en),
      .clk(clk),
      .out(mul_reg_out),
      .done(mul_reg_done)
  );
  
  std_reg #(32) acc (
      .in(acc_in),
      .write_en(acc_write_en),
      .clk(clk),
      .out(acc_out),
      .done(acc_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign down = top;
  assign right = left;
  assign out = acc_out;
  assign done = (fsm0_out == 32'd2) ? 1'd1 : '0;
  assign mul_left = (fsm0_out == 32'd0 & !mul_reg_done & go) ? top : '0;
  assign mul_right = (fsm0_out == 32'd0 & !mul_reg_done & go) ? left : '0;
  assign mul_go = (!mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign add_left = (fsm0_out == 32'd1 & !acc_done & go) ? acc_out : '0;
  assign add_right = (fsm0_out == 32'd1 & !acc_done & go) ? mul_reg_out : '0;
  assign mul_reg_in = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? mul_out : '0;
  assign mul_reg_write_en = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign acc_in = (fsm0_out == 32'd1 & !acc_done & go) ? add_out : '0;
  assign acc_write_en = (fsm0_out == 32'd1 & !acc_done & go) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd1 & acc_done & go) ? 32'd2 : (fsm0_out == 32'd0 & mul_reg_done & go) ? 32'd1 : (fsm0_out == 32'd2) ? 32'd0 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & mul_reg_done & go | fsm0_out == 32'd1 & acc_done & go | fsm0_out == 32'd2) ? 1'd1 : '0;
endmodule // end mac_pe
// Component Signature
module main (
      input wire go,
      input wire clk,
      input wire [31:0] out_mem_read_data,
      input wire out_mem_done,
      output wire done,
      output wire [2:0] out_mem_addr0,
      output wire [2:0] out_mem_addr1,
      output wire [31:0] out_mem_write_data,
      output wire out_mem_write_en
  );
  
  // Structure wire declarations
  wire [31:0] left_44_read_in;
  wire left_44_read_write_en;
  wire left_44_read_clk;
  wire [31:0] left_44_read_out;
  wire left_44_read_done;
  wire [31:0] top_44_read_in;
  wire top_44_read_write_en;
  wire top_44_read_clk;
  wire [31:0] top_44_read_out;
  wire top_44_read_done;
  wire [31:0] pe_44_top;
  wire [31:0] pe_44_left;
  wire pe_44_go;
  wire pe_44_clk;
  wire [31:0] pe_44_down;
  wire [31:0] pe_44_right;
  wire [31:0] pe_44_out;
  wire pe_44_done;
  wire [31:0] right_43_write_in;
  wire right_43_write_write_en;
  wire right_43_write_clk;
  wire [31:0] right_43_write_out;
  wire right_43_write_done;
  wire [31:0] left_43_read_in;
  wire left_43_read_write_en;
  wire left_43_read_clk;
  wire [31:0] left_43_read_out;
  wire left_43_read_done;
  wire [31:0] top_43_read_in;
  wire top_43_read_write_en;
  wire top_43_read_clk;
  wire [31:0] top_43_read_out;
  wire top_43_read_done;
  wire [31:0] pe_43_top;
  wire [31:0] pe_43_left;
  wire pe_43_go;
  wire pe_43_clk;
  wire [31:0] pe_43_down;
  wire [31:0] pe_43_right;
  wire [31:0] pe_43_out;
  wire pe_43_done;
  wire [31:0] right_42_write_in;
  wire right_42_write_write_en;
  wire right_42_write_clk;
  wire [31:0] right_42_write_out;
  wire right_42_write_done;
  wire [31:0] left_42_read_in;
  wire left_42_read_write_en;
  wire left_42_read_clk;
  wire [31:0] left_42_read_out;
  wire left_42_read_done;
  wire [31:0] top_42_read_in;
  wire top_42_read_write_en;
  wire top_42_read_clk;
  wire [31:0] top_42_read_out;
  wire top_42_read_done;
  wire [31:0] pe_42_top;
  wire [31:0] pe_42_left;
  wire pe_42_go;
  wire pe_42_clk;
  wire [31:0] pe_42_down;
  wire [31:0] pe_42_right;
  wire [31:0] pe_42_out;
  wire pe_42_done;
  wire [31:0] right_41_write_in;
  wire right_41_write_write_en;
  wire right_41_write_clk;
  wire [31:0] right_41_write_out;
  wire right_41_write_done;
  wire [31:0] left_41_read_in;
  wire left_41_read_write_en;
  wire left_41_read_clk;
  wire [31:0] left_41_read_out;
  wire left_41_read_done;
  wire [31:0] top_41_read_in;
  wire top_41_read_write_en;
  wire top_41_read_clk;
  wire [31:0] top_41_read_out;
  wire top_41_read_done;
  wire [31:0] pe_41_top;
  wire [31:0] pe_41_left;
  wire pe_41_go;
  wire pe_41_clk;
  wire [31:0] pe_41_down;
  wire [31:0] pe_41_right;
  wire [31:0] pe_41_out;
  wire pe_41_done;
  wire [31:0] right_40_write_in;
  wire right_40_write_write_en;
  wire right_40_write_clk;
  wire [31:0] right_40_write_out;
  wire right_40_write_done;
  wire [31:0] left_40_read_in;
  wire left_40_read_write_en;
  wire left_40_read_clk;
  wire [31:0] left_40_read_out;
  wire left_40_read_done;
  wire [31:0] top_40_read_in;
  wire top_40_read_write_en;
  wire top_40_read_clk;
  wire [31:0] top_40_read_out;
  wire top_40_read_done;
  wire [31:0] pe_40_top;
  wire [31:0] pe_40_left;
  wire pe_40_go;
  wire pe_40_clk;
  wire [31:0] pe_40_down;
  wire [31:0] pe_40_right;
  wire [31:0] pe_40_out;
  wire pe_40_done;
  wire [31:0] down_34_write_in;
  wire down_34_write_write_en;
  wire down_34_write_clk;
  wire [31:0] down_34_write_out;
  wire down_34_write_done;
  wire [31:0] left_34_read_in;
  wire left_34_read_write_en;
  wire left_34_read_clk;
  wire [31:0] left_34_read_out;
  wire left_34_read_done;
  wire [31:0] top_34_read_in;
  wire top_34_read_write_en;
  wire top_34_read_clk;
  wire [31:0] top_34_read_out;
  wire top_34_read_done;
  wire [31:0] pe_34_top;
  wire [31:0] pe_34_left;
  wire pe_34_go;
  wire pe_34_clk;
  wire [31:0] pe_34_down;
  wire [31:0] pe_34_right;
  wire [31:0] pe_34_out;
  wire pe_34_done;
  wire [31:0] down_33_write_in;
  wire down_33_write_write_en;
  wire down_33_write_clk;
  wire [31:0] down_33_write_out;
  wire down_33_write_done;
  wire [31:0] right_33_write_in;
  wire right_33_write_write_en;
  wire right_33_write_clk;
  wire [31:0] right_33_write_out;
  wire right_33_write_done;
  wire [31:0] left_33_read_in;
  wire left_33_read_write_en;
  wire left_33_read_clk;
  wire [31:0] left_33_read_out;
  wire left_33_read_done;
  wire [31:0] top_33_read_in;
  wire top_33_read_write_en;
  wire top_33_read_clk;
  wire [31:0] top_33_read_out;
  wire top_33_read_done;
  wire [31:0] pe_33_top;
  wire [31:0] pe_33_left;
  wire pe_33_go;
  wire pe_33_clk;
  wire [31:0] pe_33_down;
  wire [31:0] pe_33_right;
  wire [31:0] pe_33_out;
  wire pe_33_done;
  wire [31:0] down_32_write_in;
  wire down_32_write_write_en;
  wire down_32_write_clk;
  wire [31:0] down_32_write_out;
  wire down_32_write_done;
  wire [31:0] right_32_write_in;
  wire right_32_write_write_en;
  wire right_32_write_clk;
  wire [31:0] right_32_write_out;
  wire right_32_write_done;
  wire [31:0] left_32_read_in;
  wire left_32_read_write_en;
  wire left_32_read_clk;
  wire [31:0] left_32_read_out;
  wire left_32_read_done;
  wire [31:0] top_32_read_in;
  wire top_32_read_write_en;
  wire top_32_read_clk;
  wire [31:0] top_32_read_out;
  wire top_32_read_done;
  wire [31:0] pe_32_top;
  wire [31:0] pe_32_left;
  wire pe_32_go;
  wire pe_32_clk;
  wire [31:0] pe_32_down;
  wire [31:0] pe_32_right;
  wire [31:0] pe_32_out;
  wire pe_32_done;
  wire [31:0] down_31_write_in;
  wire down_31_write_write_en;
  wire down_31_write_clk;
  wire [31:0] down_31_write_out;
  wire down_31_write_done;
  wire [31:0] right_31_write_in;
  wire right_31_write_write_en;
  wire right_31_write_clk;
  wire [31:0] right_31_write_out;
  wire right_31_write_done;
  wire [31:0] left_31_read_in;
  wire left_31_read_write_en;
  wire left_31_read_clk;
  wire [31:0] left_31_read_out;
  wire left_31_read_done;
  wire [31:0] top_31_read_in;
  wire top_31_read_write_en;
  wire top_31_read_clk;
  wire [31:0] top_31_read_out;
  wire top_31_read_done;
  wire [31:0] pe_31_top;
  wire [31:0] pe_31_left;
  wire pe_31_go;
  wire pe_31_clk;
  wire [31:0] pe_31_down;
  wire [31:0] pe_31_right;
  wire [31:0] pe_31_out;
  wire pe_31_done;
  wire [31:0] down_30_write_in;
  wire down_30_write_write_en;
  wire down_30_write_clk;
  wire [31:0] down_30_write_out;
  wire down_30_write_done;
  wire [31:0] right_30_write_in;
  wire right_30_write_write_en;
  wire right_30_write_clk;
  wire [31:0] right_30_write_out;
  wire right_30_write_done;
  wire [31:0] left_30_read_in;
  wire left_30_read_write_en;
  wire left_30_read_clk;
  wire [31:0] left_30_read_out;
  wire left_30_read_done;
  wire [31:0] top_30_read_in;
  wire top_30_read_write_en;
  wire top_30_read_clk;
  wire [31:0] top_30_read_out;
  wire top_30_read_done;
  wire [31:0] pe_30_top;
  wire [31:0] pe_30_left;
  wire pe_30_go;
  wire pe_30_clk;
  wire [31:0] pe_30_down;
  wire [31:0] pe_30_right;
  wire [31:0] pe_30_out;
  wire pe_30_done;
  wire [31:0] down_24_write_in;
  wire down_24_write_write_en;
  wire down_24_write_clk;
  wire [31:0] down_24_write_out;
  wire down_24_write_done;
  wire [31:0] left_24_read_in;
  wire left_24_read_write_en;
  wire left_24_read_clk;
  wire [31:0] left_24_read_out;
  wire left_24_read_done;
  wire [31:0] top_24_read_in;
  wire top_24_read_write_en;
  wire top_24_read_clk;
  wire [31:0] top_24_read_out;
  wire top_24_read_done;
  wire [31:0] pe_24_top;
  wire [31:0] pe_24_left;
  wire pe_24_go;
  wire pe_24_clk;
  wire [31:0] pe_24_down;
  wire [31:0] pe_24_right;
  wire [31:0] pe_24_out;
  wire pe_24_done;
  wire [31:0] down_23_write_in;
  wire down_23_write_write_en;
  wire down_23_write_clk;
  wire [31:0] down_23_write_out;
  wire down_23_write_done;
  wire [31:0] right_23_write_in;
  wire right_23_write_write_en;
  wire right_23_write_clk;
  wire [31:0] right_23_write_out;
  wire right_23_write_done;
  wire [31:0] left_23_read_in;
  wire left_23_read_write_en;
  wire left_23_read_clk;
  wire [31:0] left_23_read_out;
  wire left_23_read_done;
  wire [31:0] top_23_read_in;
  wire top_23_read_write_en;
  wire top_23_read_clk;
  wire [31:0] top_23_read_out;
  wire top_23_read_done;
  wire [31:0] pe_23_top;
  wire [31:0] pe_23_left;
  wire pe_23_go;
  wire pe_23_clk;
  wire [31:0] pe_23_down;
  wire [31:0] pe_23_right;
  wire [31:0] pe_23_out;
  wire pe_23_done;
  wire [31:0] down_22_write_in;
  wire down_22_write_write_en;
  wire down_22_write_clk;
  wire [31:0] down_22_write_out;
  wire down_22_write_done;
  wire [31:0] right_22_write_in;
  wire right_22_write_write_en;
  wire right_22_write_clk;
  wire [31:0] right_22_write_out;
  wire right_22_write_done;
  wire [31:0] left_22_read_in;
  wire left_22_read_write_en;
  wire left_22_read_clk;
  wire [31:0] left_22_read_out;
  wire left_22_read_done;
  wire [31:0] top_22_read_in;
  wire top_22_read_write_en;
  wire top_22_read_clk;
  wire [31:0] top_22_read_out;
  wire top_22_read_done;
  wire [31:0] pe_22_top;
  wire [31:0] pe_22_left;
  wire pe_22_go;
  wire pe_22_clk;
  wire [31:0] pe_22_down;
  wire [31:0] pe_22_right;
  wire [31:0] pe_22_out;
  wire pe_22_done;
  wire [31:0] down_21_write_in;
  wire down_21_write_write_en;
  wire down_21_write_clk;
  wire [31:0] down_21_write_out;
  wire down_21_write_done;
  wire [31:0] right_21_write_in;
  wire right_21_write_write_en;
  wire right_21_write_clk;
  wire [31:0] right_21_write_out;
  wire right_21_write_done;
  wire [31:0] left_21_read_in;
  wire left_21_read_write_en;
  wire left_21_read_clk;
  wire [31:0] left_21_read_out;
  wire left_21_read_done;
  wire [31:0] top_21_read_in;
  wire top_21_read_write_en;
  wire top_21_read_clk;
  wire [31:0] top_21_read_out;
  wire top_21_read_done;
  wire [31:0] pe_21_top;
  wire [31:0] pe_21_left;
  wire pe_21_go;
  wire pe_21_clk;
  wire [31:0] pe_21_down;
  wire [31:0] pe_21_right;
  wire [31:0] pe_21_out;
  wire pe_21_done;
  wire [31:0] down_20_write_in;
  wire down_20_write_write_en;
  wire down_20_write_clk;
  wire [31:0] down_20_write_out;
  wire down_20_write_done;
  wire [31:0] right_20_write_in;
  wire right_20_write_write_en;
  wire right_20_write_clk;
  wire [31:0] right_20_write_out;
  wire right_20_write_done;
  wire [31:0] left_20_read_in;
  wire left_20_read_write_en;
  wire left_20_read_clk;
  wire [31:0] left_20_read_out;
  wire left_20_read_done;
  wire [31:0] top_20_read_in;
  wire top_20_read_write_en;
  wire top_20_read_clk;
  wire [31:0] top_20_read_out;
  wire top_20_read_done;
  wire [31:0] pe_20_top;
  wire [31:0] pe_20_left;
  wire pe_20_go;
  wire pe_20_clk;
  wire [31:0] pe_20_down;
  wire [31:0] pe_20_right;
  wire [31:0] pe_20_out;
  wire pe_20_done;
  wire [31:0] down_14_write_in;
  wire down_14_write_write_en;
  wire down_14_write_clk;
  wire [31:0] down_14_write_out;
  wire down_14_write_done;
  wire [31:0] left_14_read_in;
  wire left_14_read_write_en;
  wire left_14_read_clk;
  wire [31:0] left_14_read_out;
  wire left_14_read_done;
  wire [31:0] top_14_read_in;
  wire top_14_read_write_en;
  wire top_14_read_clk;
  wire [31:0] top_14_read_out;
  wire top_14_read_done;
  wire [31:0] pe_14_top;
  wire [31:0] pe_14_left;
  wire pe_14_go;
  wire pe_14_clk;
  wire [31:0] pe_14_down;
  wire [31:0] pe_14_right;
  wire [31:0] pe_14_out;
  wire pe_14_done;
  wire [31:0] down_13_write_in;
  wire down_13_write_write_en;
  wire down_13_write_clk;
  wire [31:0] down_13_write_out;
  wire down_13_write_done;
  wire [31:0] right_13_write_in;
  wire right_13_write_write_en;
  wire right_13_write_clk;
  wire [31:0] right_13_write_out;
  wire right_13_write_done;
  wire [31:0] left_13_read_in;
  wire left_13_read_write_en;
  wire left_13_read_clk;
  wire [31:0] left_13_read_out;
  wire left_13_read_done;
  wire [31:0] top_13_read_in;
  wire top_13_read_write_en;
  wire top_13_read_clk;
  wire [31:0] top_13_read_out;
  wire top_13_read_done;
  wire [31:0] pe_13_top;
  wire [31:0] pe_13_left;
  wire pe_13_go;
  wire pe_13_clk;
  wire [31:0] pe_13_down;
  wire [31:0] pe_13_right;
  wire [31:0] pe_13_out;
  wire pe_13_done;
  wire [31:0] down_12_write_in;
  wire down_12_write_write_en;
  wire down_12_write_clk;
  wire [31:0] down_12_write_out;
  wire down_12_write_done;
  wire [31:0] right_12_write_in;
  wire right_12_write_write_en;
  wire right_12_write_clk;
  wire [31:0] right_12_write_out;
  wire right_12_write_done;
  wire [31:0] left_12_read_in;
  wire left_12_read_write_en;
  wire left_12_read_clk;
  wire [31:0] left_12_read_out;
  wire left_12_read_done;
  wire [31:0] top_12_read_in;
  wire top_12_read_write_en;
  wire top_12_read_clk;
  wire [31:0] top_12_read_out;
  wire top_12_read_done;
  wire [31:0] pe_12_top;
  wire [31:0] pe_12_left;
  wire pe_12_go;
  wire pe_12_clk;
  wire [31:0] pe_12_down;
  wire [31:0] pe_12_right;
  wire [31:0] pe_12_out;
  wire pe_12_done;
  wire [31:0] down_11_write_in;
  wire down_11_write_write_en;
  wire down_11_write_clk;
  wire [31:0] down_11_write_out;
  wire down_11_write_done;
  wire [31:0] right_11_write_in;
  wire right_11_write_write_en;
  wire right_11_write_clk;
  wire [31:0] right_11_write_out;
  wire right_11_write_done;
  wire [31:0] left_11_read_in;
  wire left_11_read_write_en;
  wire left_11_read_clk;
  wire [31:0] left_11_read_out;
  wire left_11_read_done;
  wire [31:0] top_11_read_in;
  wire top_11_read_write_en;
  wire top_11_read_clk;
  wire [31:0] top_11_read_out;
  wire top_11_read_done;
  wire [31:0] pe_11_top;
  wire [31:0] pe_11_left;
  wire pe_11_go;
  wire pe_11_clk;
  wire [31:0] pe_11_down;
  wire [31:0] pe_11_right;
  wire [31:0] pe_11_out;
  wire pe_11_done;
  wire [31:0] down_10_write_in;
  wire down_10_write_write_en;
  wire down_10_write_clk;
  wire [31:0] down_10_write_out;
  wire down_10_write_done;
  wire [31:0] right_10_write_in;
  wire right_10_write_write_en;
  wire right_10_write_clk;
  wire [31:0] right_10_write_out;
  wire right_10_write_done;
  wire [31:0] left_10_read_in;
  wire left_10_read_write_en;
  wire left_10_read_clk;
  wire [31:0] left_10_read_out;
  wire left_10_read_done;
  wire [31:0] top_10_read_in;
  wire top_10_read_write_en;
  wire top_10_read_clk;
  wire [31:0] top_10_read_out;
  wire top_10_read_done;
  wire [31:0] pe_10_top;
  wire [31:0] pe_10_left;
  wire pe_10_go;
  wire pe_10_clk;
  wire [31:0] pe_10_down;
  wire [31:0] pe_10_right;
  wire [31:0] pe_10_out;
  wire pe_10_done;
  wire [31:0] down_04_write_in;
  wire down_04_write_write_en;
  wire down_04_write_clk;
  wire [31:0] down_04_write_out;
  wire down_04_write_done;
  wire [31:0] left_04_read_in;
  wire left_04_read_write_en;
  wire left_04_read_clk;
  wire [31:0] left_04_read_out;
  wire left_04_read_done;
  wire [31:0] top_04_read_in;
  wire top_04_read_write_en;
  wire top_04_read_clk;
  wire [31:0] top_04_read_out;
  wire top_04_read_done;
  wire [31:0] pe_04_top;
  wire [31:0] pe_04_left;
  wire pe_04_go;
  wire pe_04_clk;
  wire [31:0] pe_04_down;
  wire [31:0] pe_04_right;
  wire [31:0] pe_04_out;
  wire pe_04_done;
  wire [31:0] down_03_write_in;
  wire down_03_write_write_en;
  wire down_03_write_clk;
  wire [31:0] down_03_write_out;
  wire down_03_write_done;
  wire [31:0] right_03_write_in;
  wire right_03_write_write_en;
  wire right_03_write_clk;
  wire [31:0] right_03_write_out;
  wire right_03_write_done;
  wire [31:0] left_03_read_in;
  wire left_03_read_write_en;
  wire left_03_read_clk;
  wire [31:0] left_03_read_out;
  wire left_03_read_done;
  wire [31:0] top_03_read_in;
  wire top_03_read_write_en;
  wire top_03_read_clk;
  wire [31:0] top_03_read_out;
  wire top_03_read_done;
  wire [31:0] pe_03_top;
  wire [31:0] pe_03_left;
  wire pe_03_go;
  wire pe_03_clk;
  wire [31:0] pe_03_down;
  wire [31:0] pe_03_right;
  wire [31:0] pe_03_out;
  wire pe_03_done;
  wire [31:0] down_02_write_in;
  wire down_02_write_write_en;
  wire down_02_write_clk;
  wire [31:0] down_02_write_out;
  wire down_02_write_done;
  wire [31:0] right_02_write_in;
  wire right_02_write_write_en;
  wire right_02_write_clk;
  wire [31:0] right_02_write_out;
  wire right_02_write_done;
  wire [31:0] left_02_read_in;
  wire left_02_read_write_en;
  wire left_02_read_clk;
  wire [31:0] left_02_read_out;
  wire left_02_read_done;
  wire [31:0] top_02_read_in;
  wire top_02_read_write_en;
  wire top_02_read_clk;
  wire [31:0] top_02_read_out;
  wire top_02_read_done;
  wire [31:0] pe_02_top;
  wire [31:0] pe_02_left;
  wire pe_02_go;
  wire pe_02_clk;
  wire [31:0] pe_02_down;
  wire [31:0] pe_02_right;
  wire [31:0] pe_02_out;
  wire pe_02_done;
  wire [31:0] down_01_write_in;
  wire down_01_write_write_en;
  wire down_01_write_clk;
  wire [31:0] down_01_write_out;
  wire down_01_write_done;
  wire [31:0] right_01_write_in;
  wire right_01_write_write_en;
  wire right_01_write_clk;
  wire [31:0] right_01_write_out;
  wire right_01_write_done;
  wire [31:0] left_01_read_in;
  wire left_01_read_write_en;
  wire left_01_read_clk;
  wire [31:0] left_01_read_out;
  wire left_01_read_done;
  wire [31:0] top_01_read_in;
  wire top_01_read_write_en;
  wire top_01_read_clk;
  wire [31:0] top_01_read_out;
  wire top_01_read_done;
  wire [31:0] pe_01_top;
  wire [31:0] pe_01_left;
  wire pe_01_go;
  wire pe_01_clk;
  wire [31:0] pe_01_down;
  wire [31:0] pe_01_right;
  wire [31:0] pe_01_out;
  wire pe_01_done;
  wire [31:0] down_00_write_in;
  wire down_00_write_write_en;
  wire down_00_write_clk;
  wire [31:0] down_00_write_out;
  wire down_00_write_done;
  wire [31:0] right_00_write_in;
  wire right_00_write_write_en;
  wire right_00_write_clk;
  wire [31:0] right_00_write_out;
  wire right_00_write_done;
  wire [31:0] left_00_read_in;
  wire left_00_read_write_en;
  wire left_00_read_clk;
  wire [31:0] left_00_read_out;
  wire left_00_read_done;
  wire [31:0] top_00_read_in;
  wire top_00_read_write_en;
  wire top_00_read_clk;
  wire [31:0] top_00_read_out;
  wire top_00_read_done;
  wire [31:0] pe_00_top;
  wire [31:0] pe_00_left;
  wire pe_00_go;
  wire pe_00_clk;
  wire [31:0] pe_00_down;
  wire [31:0] pe_00_right;
  wire [31:0] pe_00_out;
  wire pe_00_done;
  wire [2:0] l4_addr0;
  wire [31:0] l4_write_data;
  wire l4_write_en;
  wire l4_clk;
  wire [31:0] l4_read_data;
  wire l4_done;
  wire [2:0] l4_add_left;
  wire [2:0] l4_add_right;
  wire [2:0] l4_add_out;
  wire [2:0] l4_idx_in;
  wire l4_idx_write_en;
  wire l4_idx_clk;
  wire [2:0] l4_idx_out;
  wire l4_idx_done;
  wire [2:0] l3_addr0;
  wire [31:0] l3_write_data;
  wire l3_write_en;
  wire l3_clk;
  wire [31:0] l3_read_data;
  wire l3_done;
  wire [2:0] l3_add_left;
  wire [2:0] l3_add_right;
  wire [2:0] l3_add_out;
  wire [2:0] l3_idx_in;
  wire l3_idx_write_en;
  wire l3_idx_clk;
  wire [2:0] l3_idx_out;
  wire l3_idx_done;
  wire [2:0] l2_addr0;
  wire [31:0] l2_write_data;
  wire l2_write_en;
  wire l2_clk;
  wire [31:0] l2_read_data;
  wire l2_done;
  wire [2:0] l2_add_left;
  wire [2:0] l2_add_right;
  wire [2:0] l2_add_out;
  wire [2:0] l2_idx_in;
  wire l2_idx_write_en;
  wire l2_idx_clk;
  wire [2:0] l2_idx_out;
  wire l2_idx_done;
  wire [2:0] l1_addr0;
  wire [31:0] l1_write_data;
  wire l1_write_en;
  wire l1_clk;
  wire [31:0] l1_read_data;
  wire l1_done;
  wire [2:0] l1_add_left;
  wire [2:0] l1_add_right;
  wire [2:0] l1_add_out;
  wire [2:0] l1_idx_in;
  wire l1_idx_write_en;
  wire l1_idx_clk;
  wire [2:0] l1_idx_out;
  wire l1_idx_done;
  wire [2:0] l0_addr0;
  wire [31:0] l0_write_data;
  wire l0_write_en;
  wire l0_clk;
  wire [31:0] l0_read_data;
  wire l0_done;
  wire [2:0] l0_add_left;
  wire [2:0] l0_add_right;
  wire [2:0] l0_add_out;
  wire [2:0] l0_idx_in;
  wire l0_idx_write_en;
  wire l0_idx_clk;
  wire [2:0] l0_idx_out;
  wire l0_idx_done;
  wire [2:0] t4_addr0;
  wire [31:0] t4_write_data;
  wire t4_write_en;
  wire t4_clk;
  wire [31:0] t4_read_data;
  wire t4_done;
  wire [2:0] t4_add_left;
  wire [2:0] t4_add_right;
  wire [2:0] t4_add_out;
  wire [2:0] t4_idx_in;
  wire t4_idx_write_en;
  wire t4_idx_clk;
  wire [2:0] t4_idx_out;
  wire t4_idx_done;
  wire [2:0] t3_addr0;
  wire [31:0] t3_write_data;
  wire t3_write_en;
  wire t3_clk;
  wire [31:0] t3_read_data;
  wire t3_done;
  wire [2:0] t3_add_left;
  wire [2:0] t3_add_right;
  wire [2:0] t3_add_out;
  wire [2:0] t3_idx_in;
  wire t3_idx_write_en;
  wire t3_idx_clk;
  wire [2:0] t3_idx_out;
  wire t3_idx_done;
  wire [2:0] t2_addr0;
  wire [31:0] t2_write_data;
  wire t2_write_en;
  wire t2_clk;
  wire [31:0] t2_read_data;
  wire t2_done;
  wire [2:0] t2_add_left;
  wire [2:0] t2_add_right;
  wire [2:0] t2_add_out;
  wire [2:0] t2_idx_in;
  wire t2_idx_write_en;
  wire t2_idx_clk;
  wire [2:0] t2_idx_out;
  wire t2_idx_done;
  wire [2:0] t1_addr0;
  wire [31:0] t1_write_data;
  wire t1_write_en;
  wire t1_clk;
  wire [31:0] t1_read_data;
  wire t1_done;
  wire [2:0] t1_add_left;
  wire [2:0] t1_add_right;
  wire [2:0] t1_add_out;
  wire [2:0] t1_idx_in;
  wire t1_idx_write_en;
  wire t1_idx_clk;
  wire [2:0] t1_idx_out;
  wire t1_idx_done;
  wire [2:0] t0_addr0;
  wire [31:0] t0_write_data;
  wire t0_write_en;
  wire t0_clk;
  wire [31:0] t0_read_data;
  wire t0_done;
  wire [2:0] t0_add_left;
  wire [2:0] t0_add_right;
  wire [2:0] t0_add_out;
  wire [2:0] t0_idx_in;
  wire t0_idx_write_en;
  wire t0_idx_clk;
  wire [2:0] t0_idx_out;
  wire t0_idx_done;
  wire par_reset0_in;
  wire par_reset0_write_en;
  wire par_reset0_clk;
  wire par_reset0_out;
  wire par_reset0_done;
  wire par_done_reg0_in;
  wire par_done_reg0_write_en;
  wire par_done_reg0_clk;
  wire par_done_reg0_out;
  wire par_done_reg0_done;
  wire par_done_reg1_in;
  wire par_done_reg1_write_en;
  wire par_done_reg1_clk;
  wire par_done_reg1_out;
  wire par_done_reg1_done;
  wire par_done_reg2_in;
  wire par_done_reg2_write_en;
  wire par_done_reg2_clk;
  wire par_done_reg2_out;
  wire par_done_reg2_done;
  wire par_done_reg3_in;
  wire par_done_reg3_write_en;
  wire par_done_reg3_clk;
  wire par_done_reg3_out;
  wire par_done_reg3_done;
  wire par_done_reg4_in;
  wire par_done_reg4_write_en;
  wire par_done_reg4_clk;
  wire par_done_reg4_out;
  wire par_done_reg4_done;
  wire par_done_reg5_in;
  wire par_done_reg5_write_en;
  wire par_done_reg5_clk;
  wire par_done_reg5_out;
  wire par_done_reg5_done;
  wire par_done_reg6_in;
  wire par_done_reg6_write_en;
  wire par_done_reg6_clk;
  wire par_done_reg6_out;
  wire par_done_reg6_done;
  wire par_done_reg7_in;
  wire par_done_reg7_write_en;
  wire par_done_reg7_clk;
  wire par_done_reg7_out;
  wire par_done_reg7_done;
  wire par_done_reg8_in;
  wire par_done_reg8_write_en;
  wire par_done_reg8_clk;
  wire par_done_reg8_out;
  wire par_done_reg8_done;
  wire par_done_reg9_in;
  wire par_done_reg9_write_en;
  wire par_done_reg9_clk;
  wire par_done_reg9_out;
  wire par_done_reg9_done;
  wire par_reset1_in;
  wire par_reset1_write_en;
  wire par_reset1_clk;
  wire par_reset1_out;
  wire par_reset1_done;
  wire par_done_reg10_in;
  wire par_done_reg10_write_en;
  wire par_done_reg10_clk;
  wire par_done_reg10_out;
  wire par_done_reg10_done;
  wire par_done_reg11_in;
  wire par_done_reg11_write_en;
  wire par_done_reg11_clk;
  wire par_done_reg11_out;
  wire par_done_reg11_done;
  wire par_reset2_in;
  wire par_reset2_write_en;
  wire par_reset2_clk;
  wire par_reset2_out;
  wire par_reset2_done;
  wire par_done_reg12_in;
  wire par_done_reg12_write_en;
  wire par_done_reg12_clk;
  wire par_done_reg12_out;
  wire par_done_reg12_done;
  wire par_done_reg13_in;
  wire par_done_reg13_write_en;
  wire par_done_reg13_clk;
  wire par_done_reg13_out;
  wire par_done_reg13_done;
  wire par_reset3_in;
  wire par_reset3_write_en;
  wire par_reset3_clk;
  wire par_reset3_out;
  wire par_reset3_done;
  wire par_done_reg14_in;
  wire par_done_reg14_write_en;
  wire par_done_reg14_clk;
  wire par_done_reg14_out;
  wire par_done_reg14_done;
  wire par_done_reg15_in;
  wire par_done_reg15_write_en;
  wire par_done_reg15_clk;
  wire par_done_reg15_out;
  wire par_done_reg15_done;
  wire par_done_reg16_in;
  wire par_done_reg16_write_en;
  wire par_done_reg16_clk;
  wire par_done_reg16_out;
  wire par_done_reg16_done;
  wire par_done_reg17_in;
  wire par_done_reg17_write_en;
  wire par_done_reg17_clk;
  wire par_done_reg17_out;
  wire par_done_reg17_done;
  wire par_done_reg18_in;
  wire par_done_reg18_write_en;
  wire par_done_reg18_clk;
  wire par_done_reg18_out;
  wire par_done_reg18_done;
  wire par_reset4_in;
  wire par_reset4_write_en;
  wire par_reset4_clk;
  wire par_reset4_out;
  wire par_reset4_done;
  wire par_done_reg19_in;
  wire par_done_reg19_write_en;
  wire par_done_reg19_clk;
  wire par_done_reg19_out;
  wire par_done_reg19_done;
  wire par_done_reg20_in;
  wire par_done_reg20_write_en;
  wire par_done_reg20_clk;
  wire par_done_reg20_out;
  wire par_done_reg20_done;
  wire par_done_reg21_in;
  wire par_done_reg21_write_en;
  wire par_done_reg21_clk;
  wire par_done_reg21_out;
  wire par_done_reg21_done;
  wire par_done_reg22_in;
  wire par_done_reg22_write_en;
  wire par_done_reg22_clk;
  wire par_done_reg22_out;
  wire par_done_reg22_done;
  wire par_done_reg23_in;
  wire par_done_reg23_write_en;
  wire par_done_reg23_clk;
  wire par_done_reg23_out;
  wire par_done_reg23_done;
  wire par_done_reg24_in;
  wire par_done_reg24_write_en;
  wire par_done_reg24_clk;
  wire par_done_reg24_out;
  wire par_done_reg24_done;
  wire par_reset5_in;
  wire par_reset5_write_en;
  wire par_reset5_clk;
  wire par_reset5_out;
  wire par_reset5_done;
  wire par_done_reg25_in;
  wire par_done_reg25_write_en;
  wire par_done_reg25_clk;
  wire par_done_reg25_out;
  wire par_done_reg25_done;
  wire par_done_reg26_in;
  wire par_done_reg26_write_en;
  wire par_done_reg26_clk;
  wire par_done_reg26_out;
  wire par_done_reg26_done;
  wire par_done_reg27_in;
  wire par_done_reg27_write_en;
  wire par_done_reg27_clk;
  wire par_done_reg27_out;
  wire par_done_reg27_done;
  wire par_done_reg28_in;
  wire par_done_reg28_write_en;
  wire par_done_reg28_clk;
  wire par_done_reg28_out;
  wire par_done_reg28_done;
  wire par_done_reg29_in;
  wire par_done_reg29_write_en;
  wire par_done_reg29_clk;
  wire par_done_reg29_out;
  wire par_done_reg29_done;
  wire par_done_reg30_in;
  wire par_done_reg30_write_en;
  wire par_done_reg30_clk;
  wire par_done_reg30_out;
  wire par_done_reg30_done;
  wire par_done_reg31_in;
  wire par_done_reg31_write_en;
  wire par_done_reg31_clk;
  wire par_done_reg31_out;
  wire par_done_reg31_done;
  wire par_done_reg32_in;
  wire par_done_reg32_write_en;
  wire par_done_reg32_clk;
  wire par_done_reg32_out;
  wire par_done_reg32_done;
  wire par_done_reg33_in;
  wire par_done_reg33_write_en;
  wire par_done_reg33_clk;
  wire par_done_reg33_out;
  wire par_done_reg33_done;
  wire par_reset6_in;
  wire par_reset6_write_en;
  wire par_reset6_clk;
  wire par_reset6_out;
  wire par_reset6_done;
  wire par_done_reg34_in;
  wire par_done_reg34_write_en;
  wire par_done_reg34_clk;
  wire par_done_reg34_out;
  wire par_done_reg34_done;
  wire par_done_reg35_in;
  wire par_done_reg35_write_en;
  wire par_done_reg35_clk;
  wire par_done_reg35_out;
  wire par_done_reg35_done;
  wire par_done_reg36_in;
  wire par_done_reg36_write_en;
  wire par_done_reg36_clk;
  wire par_done_reg36_out;
  wire par_done_reg36_done;
  wire par_done_reg37_in;
  wire par_done_reg37_write_en;
  wire par_done_reg37_clk;
  wire par_done_reg37_out;
  wire par_done_reg37_done;
  wire par_done_reg38_in;
  wire par_done_reg38_write_en;
  wire par_done_reg38_clk;
  wire par_done_reg38_out;
  wire par_done_reg38_done;
  wire par_done_reg39_in;
  wire par_done_reg39_write_en;
  wire par_done_reg39_clk;
  wire par_done_reg39_out;
  wire par_done_reg39_done;
  wire par_done_reg40_in;
  wire par_done_reg40_write_en;
  wire par_done_reg40_clk;
  wire par_done_reg40_out;
  wire par_done_reg40_done;
  wire par_done_reg41_in;
  wire par_done_reg41_write_en;
  wire par_done_reg41_clk;
  wire par_done_reg41_out;
  wire par_done_reg41_done;
  wire par_done_reg42_in;
  wire par_done_reg42_write_en;
  wire par_done_reg42_clk;
  wire par_done_reg42_out;
  wire par_done_reg42_done;
  wire par_done_reg43_in;
  wire par_done_reg43_write_en;
  wire par_done_reg43_clk;
  wire par_done_reg43_out;
  wire par_done_reg43_done;
  wire par_done_reg44_in;
  wire par_done_reg44_write_en;
  wire par_done_reg44_clk;
  wire par_done_reg44_out;
  wire par_done_reg44_done;
  wire par_done_reg45_in;
  wire par_done_reg45_write_en;
  wire par_done_reg45_clk;
  wire par_done_reg45_out;
  wire par_done_reg45_done;
  wire par_reset7_in;
  wire par_reset7_write_en;
  wire par_reset7_clk;
  wire par_reset7_out;
  wire par_reset7_done;
  wire par_done_reg46_in;
  wire par_done_reg46_write_en;
  wire par_done_reg46_clk;
  wire par_done_reg46_out;
  wire par_done_reg46_done;
  wire par_done_reg47_in;
  wire par_done_reg47_write_en;
  wire par_done_reg47_clk;
  wire par_done_reg47_out;
  wire par_done_reg47_done;
  wire par_done_reg48_in;
  wire par_done_reg48_write_en;
  wire par_done_reg48_clk;
  wire par_done_reg48_out;
  wire par_done_reg48_done;
  wire par_done_reg49_in;
  wire par_done_reg49_write_en;
  wire par_done_reg49_clk;
  wire par_done_reg49_out;
  wire par_done_reg49_done;
  wire par_done_reg50_in;
  wire par_done_reg50_write_en;
  wire par_done_reg50_clk;
  wire par_done_reg50_out;
  wire par_done_reg50_done;
  wire par_done_reg51_in;
  wire par_done_reg51_write_en;
  wire par_done_reg51_clk;
  wire par_done_reg51_out;
  wire par_done_reg51_done;
  wire par_done_reg52_in;
  wire par_done_reg52_write_en;
  wire par_done_reg52_clk;
  wire par_done_reg52_out;
  wire par_done_reg52_done;
  wire par_done_reg53_in;
  wire par_done_reg53_write_en;
  wire par_done_reg53_clk;
  wire par_done_reg53_out;
  wire par_done_reg53_done;
  wire par_done_reg54_in;
  wire par_done_reg54_write_en;
  wire par_done_reg54_clk;
  wire par_done_reg54_out;
  wire par_done_reg54_done;
  wire par_done_reg55_in;
  wire par_done_reg55_write_en;
  wire par_done_reg55_clk;
  wire par_done_reg55_out;
  wire par_done_reg55_done;
  wire par_done_reg56_in;
  wire par_done_reg56_write_en;
  wire par_done_reg56_clk;
  wire par_done_reg56_out;
  wire par_done_reg56_done;
  wire par_done_reg57_in;
  wire par_done_reg57_write_en;
  wire par_done_reg57_clk;
  wire par_done_reg57_out;
  wire par_done_reg57_done;
  wire par_done_reg58_in;
  wire par_done_reg58_write_en;
  wire par_done_reg58_clk;
  wire par_done_reg58_out;
  wire par_done_reg58_done;
  wire par_done_reg59_in;
  wire par_done_reg59_write_en;
  wire par_done_reg59_clk;
  wire par_done_reg59_out;
  wire par_done_reg59_done;
  wire par_reset8_in;
  wire par_reset8_write_en;
  wire par_reset8_clk;
  wire par_reset8_out;
  wire par_reset8_done;
  wire par_done_reg60_in;
  wire par_done_reg60_write_en;
  wire par_done_reg60_clk;
  wire par_done_reg60_out;
  wire par_done_reg60_done;
  wire par_done_reg61_in;
  wire par_done_reg61_write_en;
  wire par_done_reg61_clk;
  wire par_done_reg61_out;
  wire par_done_reg61_done;
  wire par_done_reg62_in;
  wire par_done_reg62_write_en;
  wire par_done_reg62_clk;
  wire par_done_reg62_out;
  wire par_done_reg62_done;
  wire par_done_reg63_in;
  wire par_done_reg63_write_en;
  wire par_done_reg63_clk;
  wire par_done_reg63_out;
  wire par_done_reg63_done;
  wire par_done_reg64_in;
  wire par_done_reg64_write_en;
  wire par_done_reg64_clk;
  wire par_done_reg64_out;
  wire par_done_reg64_done;
  wire par_done_reg65_in;
  wire par_done_reg65_write_en;
  wire par_done_reg65_clk;
  wire par_done_reg65_out;
  wire par_done_reg65_done;
  wire par_done_reg66_in;
  wire par_done_reg66_write_en;
  wire par_done_reg66_clk;
  wire par_done_reg66_out;
  wire par_done_reg66_done;
  wire par_done_reg67_in;
  wire par_done_reg67_write_en;
  wire par_done_reg67_clk;
  wire par_done_reg67_out;
  wire par_done_reg67_done;
  wire par_done_reg68_in;
  wire par_done_reg68_write_en;
  wire par_done_reg68_clk;
  wire par_done_reg68_out;
  wire par_done_reg68_done;
  wire par_done_reg69_in;
  wire par_done_reg69_write_en;
  wire par_done_reg69_clk;
  wire par_done_reg69_out;
  wire par_done_reg69_done;
  wire par_done_reg70_in;
  wire par_done_reg70_write_en;
  wire par_done_reg70_clk;
  wire par_done_reg70_out;
  wire par_done_reg70_done;
  wire par_done_reg71_in;
  wire par_done_reg71_write_en;
  wire par_done_reg71_clk;
  wire par_done_reg71_out;
  wire par_done_reg71_done;
  wire par_done_reg72_in;
  wire par_done_reg72_write_en;
  wire par_done_reg72_clk;
  wire par_done_reg72_out;
  wire par_done_reg72_done;
  wire par_done_reg73_in;
  wire par_done_reg73_write_en;
  wire par_done_reg73_clk;
  wire par_done_reg73_out;
  wire par_done_reg73_done;
  wire par_done_reg74_in;
  wire par_done_reg74_write_en;
  wire par_done_reg74_clk;
  wire par_done_reg74_out;
  wire par_done_reg74_done;
  wire par_done_reg75_in;
  wire par_done_reg75_write_en;
  wire par_done_reg75_clk;
  wire par_done_reg75_out;
  wire par_done_reg75_done;
  wire par_done_reg76_in;
  wire par_done_reg76_write_en;
  wire par_done_reg76_clk;
  wire par_done_reg76_out;
  wire par_done_reg76_done;
  wire par_done_reg77_in;
  wire par_done_reg77_write_en;
  wire par_done_reg77_clk;
  wire par_done_reg77_out;
  wire par_done_reg77_done;
  wire par_done_reg78_in;
  wire par_done_reg78_write_en;
  wire par_done_reg78_clk;
  wire par_done_reg78_out;
  wire par_done_reg78_done;
  wire par_done_reg79_in;
  wire par_done_reg79_write_en;
  wire par_done_reg79_clk;
  wire par_done_reg79_out;
  wire par_done_reg79_done;
  wire par_reset9_in;
  wire par_reset9_write_en;
  wire par_reset9_clk;
  wire par_reset9_out;
  wire par_reset9_done;
  wire par_done_reg80_in;
  wire par_done_reg80_write_en;
  wire par_done_reg80_clk;
  wire par_done_reg80_out;
  wire par_done_reg80_done;
  wire par_done_reg81_in;
  wire par_done_reg81_write_en;
  wire par_done_reg81_clk;
  wire par_done_reg81_out;
  wire par_done_reg81_done;
  wire par_done_reg82_in;
  wire par_done_reg82_write_en;
  wire par_done_reg82_clk;
  wire par_done_reg82_out;
  wire par_done_reg82_done;
  wire par_done_reg83_in;
  wire par_done_reg83_write_en;
  wire par_done_reg83_clk;
  wire par_done_reg83_out;
  wire par_done_reg83_done;
  wire par_done_reg84_in;
  wire par_done_reg84_write_en;
  wire par_done_reg84_clk;
  wire par_done_reg84_out;
  wire par_done_reg84_done;
  wire par_done_reg85_in;
  wire par_done_reg85_write_en;
  wire par_done_reg85_clk;
  wire par_done_reg85_out;
  wire par_done_reg85_done;
  wire par_done_reg86_in;
  wire par_done_reg86_write_en;
  wire par_done_reg86_clk;
  wire par_done_reg86_out;
  wire par_done_reg86_done;
  wire par_done_reg87_in;
  wire par_done_reg87_write_en;
  wire par_done_reg87_clk;
  wire par_done_reg87_out;
  wire par_done_reg87_done;
  wire par_done_reg88_in;
  wire par_done_reg88_write_en;
  wire par_done_reg88_clk;
  wire par_done_reg88_out;
  wire par_done_reg88_done;
  wire par_done_reg89_in;
  wire par_done_reg89_write_en;
  wire par_done_reg89_clk;
  wire par_done_reg89_out;
  wire par_done_reg89_done;
  wire par_done_reg90_in;
  wire par_done_reg90_write_en;
  wire par_done_reg90_clk;
  wire par_done_reg90_out;
  wire par_done_reg90_done;
  wire par_done_reg91_in;
  wire par_done_reg91_write_en;
  wire par_done_reg91_clk;
  wire par_done_reg91_out;
  wire par_done_reg91_done;
  wire par_done_reg92_in;
  wire par_done_reg92_write_en;
  wire par_done_reg92_clk;
  wire par_done_reg92_out;
  wire par_done_reg92_done;
  wire par_done_reg93_in;
  wire par_done_reg93_write_en;
  wire par_done_reg93_clk;
  wire par_done_reg93_out;
  wire par_done_reg93_done;
  wire par_done_reg94_in;
  wire par_done_reg94_write_en;
  wire par_done_reg94_clk;
  wire par_done_reg94_out;
  wire par_done_reg94_done;
  wire par_done_reg95_in;
  wire par_done_reg95_write_en;
  wire par_done_reg95_clk;
  wire par_done_reg95_out;
  wire par_done_reg95_done;
  wire par_done_reg96_in;
  wire par_done_reg96_write_en;
  wire par_done_reg96_clk;
  wire par_done_reg96_out;
  wire par_done_reg96_done;
  wire par_done_reg97_in;
  wire par_done_reg97_write_en;
  wire par_done_reg97_clk;
  wire par_done_reg97_out;
  wire par_done_reg97_done;
  wire par_done_reg98_in;
  wire par_done_reg98_write_en;
  wire par_done_reg98_clk;
  wire par_done_reg98_out;
  wire par_done_reg98_done;
  wire par_done_reg99_in;
  wire par_done_reg99_write_en;
  wire par_done_reg99_clk;
  wire par_done_reg99_out;
  wire par_done_reg99_done;
  wire par_reset10_in;
  wire par_reset10_write_en;
  wire par_reset10_clk;
  wire par_reset10_out;
  wire par_reset10_done;
  wire par_done_reg100_in;
  wire par_done_reg100_write_en;
  wire par_done_reg100_clk;
  wire par_done_reg100_out;
  wire par_done_reg100_done;
  wire par_done_reg101_in;
  wire par_done_reg101_write_en;
  wire par_done_reg101_clk;
  wire par_done_reg101_out;
  wire par_done_reg101_done;
  wire par_done_reg102_in;
  wire par_done_reg102_write_en;
  wire par_done_reg102_clk;
  wire par_done_reg102_out;
  wire par_done_reg102_done;
  wire par_done_reg103_in;
  wire par_done_reg103_write_en;
  wire par_done_reg103_clk;
  wire par_done_reg103_out;
  wire par_done_reg103_done;
  wire par_done_reg104_in;
  wire par_done_reg104_write_en;
  wire par_done_reg104_clk;
  wire par_done_reg104_out;
  wire par_done_reg104_done;
  wire par_done_reg105_in;
  wire par_done_reg105_write_en;
  wire par_done_reg105_clk;
  wire par_done_reg105_out;
  wire par_done_reg105_done;
  wire par_done_reg106_in;
  wire par_done_reg106_write_en;
  wire par_done_reg106_clk;
  wire par_done_reg106_out;
  wire par_done_reg106_done;
  wire par_done_reg107_in;
  wire par_done_reg107_write_en;
  wire par_done_reg107_clk;
  wire par_done_reg107_out;
  wire par_done_reg107_done;
  wire par_done_reg108_in;
  wire par_done_reg108_write_en;
  wire par_done_reg108_clk;
  wire par_done_reg108_out;
  wire par_done_reg108_done;
  wire par_done_reg109_in;
  wire par_done_reg109_write_en;
  wire par_done_reg109_clk;
  wire par_done_reg109_out;
  wire par_done_reg109_done;
  wire par_done_reg110_in;
  wire par_done_reg110_write_en;
  wire par_done_reg110_clk;
  wire par_done_reg110_out;
  wire par_done_reg110_done;
  wire par_done_reg111_in;
  wire par_done_reg111_write_en;
  wire par_done_reg111_clk;
  wire par_done_reg111_out;
  wire par_done_reg111_done;
  wire par_done_reg112_in;
  wire par_done_reg112_write_en;
  wire par_done_reg112_clk;
  wire par_done_reg112_out;
  wire par_done_reg112_done;
  wire par_done_reg113_in;
  wire par_done_reg113_write_en;
  wire par_done_reg113_clk;
  wire par_done_reg113_out;
  wire par_done_reg113_done;
  wire par_done_reg114_in;
  wire par_done_reg114_write_en;
  wire par_done_reg114_clk;
  wire par_done_reg114_out;
  wire par_done_reg114_done;
  wire par_done_reg115_in;
  wire par_done_reg115_write_en;
  wire par_done_reg115_clk;
  wire par_done_reg115_out;
  wire par_done_reg115_done;
  wire par_done_reg116_in;
  wire par_done_reg116_write_en;
  wire par_done_reg116_clk;
  wire par_done_reg116_out;
  wire par_done_reg116_done;
  wire par_done_reg117_in;
  wire par_done_reg117_write_en;
  wire par_done_reg117_clk;
  wire par_done_reg117_out;
  wire par_done_reg117_done;
  wire par_done_reg118_in;
  wire par_done_reg118_write_en;
  wire par_done_reg118_clk;
  wire par_done_reg118_out;
  wire par_done_reg118_done;
  wire par_done_reg119_in;
  wire par_done_reg119_write_en;
  wire par_done_reg119_clk;
  wire par_done_reg119_out;
  wire par_done_reg119_done;
  wire par_done_reg120_in;
  wire par_done_reg120_write_en;
  wire par_done_reg120_clk;
  wire par_done_reg120_out;
  wire par_done_reg120_done;
  wire par_done_reg121_in;
  wire par_done_reg121_write_en;
  wire par_done_reg121_clk;
  wire par_done_reg121_out;
  wire par_done_reg121_done;
  wire par_done_reg122_in;
  wire par_done_reg122_write_en;
  wire par_done_reg122_clk;
  wire par_done_reg122_out;
  wire par_done_reg122_done;
  wire par_done_reg123_in;
  wire par_done_reg123_write_en;
  wire par_done_reg123_clk;
  wire par_done_reg123_out;
  wire par_done_reg123_done;
  wire par_done_reg124_in;
  wire par_done_reg124_write_en;
  wire par_done_reg124_clk;
  wire par_done_reg124_out;
  wire par_done_reg124_done;
  wire par_done_reg125_in;
  wire par_done_reg125_write_en;
  wire par_done_reg125_clk;
  wire par_done_reg125_out;
  wire par_done_reg125_done;
  wire par_done_reg126_in;
  wire par_done_reg126_write_en;
  wire par_done_reg126_clk;
  wire par_done_reg126_out;
  wire par_done_reg126_done;
  wire par_done_reg127_in;
  wire par_done_reg127_write_en;
  wire par_done_reg127_clk;
  wire par_done_reg127_out;
  wire par_done_reg127_done;
  wire par_done_reg128_in;
  wire par_done_reg128_write_en;
  wire par_done_reg128_clk;
  wire par_done_reg128_out;
  wire par_done_reg128_done;
  wire par_done_reg129_in;
  wire par_done_reg129_write_en;
  wire par_done_reg129_clk;
  wire par_done_reg129_out;
  wire par_done_reg129_done;
  wire par_reset11_in;
  wire par_reset11_write_en;
  wire par_reset11_clk;
  wire par_reset11_out;
  wire par_reset11_done;
  wire par_done_reg130_in;
  wire par_done_reg130_write_en;
  wire par_done_reg130_clk;
  wire par_done_reg130_out;
  wire par_done_reg130_done;
  wire par_done_reg131_in;
  wire par_done_reg131_write_en;
  wire par_done_reg131_clk;
  wire par_done_reg131_out;
  wire par_done_reg131_done;
  wire par_done_reg132_in;
  wire par_done_reg132_write_en;
  wire par_done_reg132_clk;
  wire par_done_reg132_out;
  wire par_done_reg132_done;
  wire par_done_reg133_in;
  wire par_done_reg133_write_en;
  wire par_done_reg133_clk;
  wire par_done_reg133_out;
  wire par_done_reg133_done;
  wire par_done_reg134_in;
  wire par_done_reg134_write_en;
  wire par_done_reg134_clk;
  wire par_done_reg134_out;
  wire par_done_reg134_done;
  wire par_done_reg135_in;
  wire par_done_reg135_write_en;
  wire par_done_reg135_clk;
  wire par_done_reg135_out;
  wire par_done_reg135_done;
  wire par_done_reg136_in;
  wire par_done_reg136_write_en;
  wire par_done_reg136_clk;
  wire par_done_reg136_out;
  wire par_done_reg136_done;
  wire par_done_reg137_in;
  wire par_done_reg137_write_en;
  wire par_done_reg137_clk;
  wire par_done_reg137_out;
  wire par_done_reg137_done;
  wire par_done_reg138_in;
  wire par_done_reg138_write_en;
  wire par_done_reg138_clk;
  wire par_done_reg138_out;
  wire par_done_reg138_done;
  wire par_done_reg139_in;
  wire par_done_reg139_write_en;
  wire par_done_reg139_clk;
  wire par_done_reg139_out;
  wire par_done_reg139_done;
  wire par_done_reg140_in;
  wire par_done_reg140_write_en;
  wire par_done_reg140_clk;
  wire par_done_reg140_out;
  wire par_done_reg140_done;
  wire par_done_reg141_in;
  wire par_done_reg141_write_en;
  wire par_done_reg141_clk;
  wire par_done_reg141_out;
  wire par_done_reg141_done;
  wire par_done_reg142_in;
  wire par_done_reg142_write_en;
  wire par_done_reg142_clk;
  wire par_done_reg142_out;
  wire par_done_reg142_done;
  wire par_done_reg143_in;
  wire par_done_reg143_write_en;
  wire par_done_reg143_clk;
  wire par_done_reg143_out;
  wire par_done_reg143_done;
  wire par_done_reg144_in;
  wire par_done_reg144_write_en;
  wire par_done_reg144_clk;
  wire par_done_reg144_out;
  wire par_done_reg144_done;
  wire par_done_reg145_in;
  wire par_done_reg145_write_en;
  wire par_done_reg145_clk;
  wire par_done_reg145_out;
  wire par_done_reg145_done;
  wire par_done_reg146_in;
  wire par_done_reg146_write_en;
  wire par_done_reg146_clk;
  wire par_done_reg146_out;
  wire par_done_reg146_done;
  wire par_done_reg147_in;
  wire par_done_reg147_write_en;
  wire par_done_reg147_clk;
  wire par_done_reg147_out;
  wire par_done_reg147_done;
  wire par_done_reg148_in;
  wire par_done_reg148_write_en;
  wire par_done_reg148_clk;
  wire par_done_reg148_out;
  wire par_done_reg148_done;
  wire par_done_reg149_in;
  wire par_done_reg149_write_en;
  wire par_done_reg149_clk;
  wire par_done_reg149_out;
  wire par_done_reg149_done;
  wire par_done_reg150_in;
  wire par_done_reg150_write_en;
  wire par_done_reg150_clk;
  wire par_done_reg150_out;
  wire par_done_reg150_done;
  wire par_done_reg151_in;
  wire par_done_reg151_write_en;
  wire par_done_reg151_clk;
  wire par_done_reg151_out;
  wire par_done_reg151_done;
  wire par_done_reg152_in;
  wire par_done_reg152_write_en;
  wire par_done_reg152_clk;
  wire par_done_reg152_out;
  wire par_done_reg152_done;
  wire par_reset12_in;
  wire par_reset12_write_en;
  wire par_reset12_clk;
  wire par_reset12_out;
  wire par_reset12_done;
  wire par_done_reg153_in;
  wire par_done_reg153_write_en;
  wire par_done_reg153_clk;
  wire par_done_reg153_out;
  wire par_done_reg153_done;
  wire par_done_reg154_in;
  wire par_done_reg154_write_en;
  wire par_done_reg154_clk;
  wire par_done_reg154_out;
  wire par_done_reg154_done;
  wire par_done_reg155_in;
  wire par_done_reg155_write_en;
  wire par_done_reg155_clk;
  wire par_done_reg155_out;
  wire par_done_reg155_done;
  wire par_done_reg156_in;
  wire par_done_reg156_write_en;
  wire par_done_reg156_clk;
  wire par_done_reg156_out;
  wire par_done_reg156_done;
  wire par_done_reg157_in;
  wire par_done_reg157_write_en;
  wire par_done_reg157_clk;
  wire par_done_reg157_out;
  wire par_done_reg157_done;
  wire par_done_reg158_in;
  wire par_done_reg158_write_en;
  wire par_done_reg158_clk;
  wire par_done_reg158_out;
  wire par_done_reg158_done;
  wire par_done_reg159_in;
  wire par_done_reg159_write_en;
  wire par_done_reg159_clk;
  wire par_done_reg159_out;
  wire par_done_reg159_done;
  wire par_done_reg160_in;
  wire par_done_reg160_write_en;
  wire par_done_reg160_clk;
  wire par_done_reg160_out;
  wire par_done_reg160_done;
  wire par_done_reg161_in;
  wire par_done_reg161_write_en;
  wire par_done_reg161_clk;
  wire par_done_reg161_out;
  wire par_done_reg161_done;
  wire par_done_reg162_in;
  wire par_done_reg162_write_en;
  wire par_done_reg162_clk;
  wire par_done_reg162_out;
  wire par_done_reg162_done;
  wire par_done_reg163_in;
  wire par_done_reg163_write_en;
  wire par_done_reg163_clk;
  wire par_done_reg163_out;
  wire par_done_reg163_done;
  wire par_done_reg164_in;
  wire par_done_reg164_write_en;
  wire par_done_reg164_clk;
  wire par_done_reg164_out;
  wire par_done_reg164_done;
  wire par_done_reg165_in;
  wire par_done_reg165_write_en;
  wire par_done_reg165_clk;
  wire par_done_reg165_out;
  wire par_done_reg165_done;
  wire par_done_reg166_in;
  wire par_done_reg166_write_en;
  wire par_done_reg166_clk;
  wire par_done_reg166_out;
  wire par_done_reg166_done;
  wire par_done_reg167_in;
  wire par_done_reg167_write_en;
  wire par_done_reg167_clk;
  wire par_done_reg167_out;
  wire par_done_reg167_done;
  wire par_done_reg168_in;
  wire par_done_reg168_write_en;
  wire par_done_reg168_clk;
  wire par_done_reg168_out;
  wire par_done_reg168_done;
  wire par_done_reg169_in;
  wire par_done_reg169_write_en;
  wire par_done_reg169_clk;
  wire par_done_reg169_out;
  wire par_done_reg169_done;
  wire par_done_reg170_in;
  wire par_done_reg170_write_en;
  wire par_done_reg170_clk;
  wire par_done_reg170_out;
  wire par_done_reg170_done;
  wire par_done_reg171_in;
  wire par_done_reg171_write_en;
  wire par_done_reg171_clk;
  wire par_done_reg171_out;
  wire par_done_reg171_done;
  wire par_done_reg172_in;
  wire par_done_reg172_write_en;
  wire par_done_reg172_clk;
  wire par_done_reg172_out;
  wire par_done_reg172_done;
  wire par_done_reg173_in;
  wire par_done_reg173_write_en;
  wire par_done_reg173_clk;
  wire par_done_reg173_out;
  wire par_done_reg173_done;
  wire par_done_reg174_in;
  wire par_done_reg174_write_en;
  wire par_done_reg174_clk;
  wire par_done_reg174_out;
  wire par_done_reg174_done;
  wire par_done_reg175_in;
  wire par_done_reg175_write_en;
  wire par_done_reg175_clk;
  wire par_done_reg175_out;
  wire par_done_reg175_done;
  wire par_done_reg176_in;
  wire par_done_reg176_write_en;
  wire par_done_reg176_clk;
  wire par_done_reg176_out;
  wire par_done_reg176_done;
  wire par_done_reg177_in;
  wire par_done_reg177_write_en;
  wire par_done_reg177_clk;
  wire par_done_reg177_out;
  wire par_done_reg177_done;
  wire par_done_reg178_in;
  wire par_done_reg178_write_en;
  wire par_done_reg178_clk;
  wire par_done_reg178_out;
  wire par_done_reg178_done;
  wire par_done_reg179_in;
  wire par_done_reg179_write_en;
  wire par_done_reg179_clk;
  wire par_done_reg179_out;
  wire par_done_reg179_done;
  wire par_done_reg180_in;
  wire par_done_reg180_write_en;
  wire par_done_reg180_clk;
  wire par_done_reg180_out;
  wire par_done_reg180_done;
  wire par_done_reg181_in;
  wire par_done_reg181_write_en;
  wire par_done_reg181_clk;
  wire par_done_reg181_out;
  wire par_done_reg181_done;
  wire par_done_reg182_in;
  wire par_done_reg182_write_en;
  wire par_done_reg182_clk;
  wire par_done_reg182_out;
  wire par_done_reg182_done;
  wire par_done_reg183_in;
  wire par_done_reg183_write_en;
  wire par_done_reg183_clk;
  wire par_done_reg183_out;
  wire par_done_reg183_done;
  wire par_done_reg184_in;
  wire par_done_reg184_write_en;
  wire par_done_reg184_clk;
  wire par_done_reg184_out;
  wire par_done_reg184_done;
  wire par_done_reg185_in;
  wire par_done_reg185_write_en;
  wire par_done_reg185_clk;
  wire par_done_reg185_out;
  wire par_done_reg185_done;
  wire par_done_reg186_in;
  wire par_done_reg186_write_en;
  wire par_done_reg186_clk;
  wire par_done_reg186_out;
  wire par_done_reg186_done;
  wire par_done_reg187_in;
  wire par_done_reg187_write_en;
  wire par_done_reg187_clk;
  wire par_done_reg187_out;
  wire par_done_reg187_done;
  wire par_done_reg188_in;
  wire par_done_reg188_write_en;
  wire par_done_reg188_clk;
  wire par_done_reg188_out;
  wire par_done_reg188_done;
  wire par_reset13_in;
  wire par_reset13_write_en;
  wire par_reset13_clk;
  wire par_reset13_out;
  wire par_reset13_done;
  wire par_done_reg189_in;
  wire par_done_reg189_write_en;
  wire par_done_reg189_clk;
  wire par_done_reg189_out;
  wire par_done_reg189_done;
  wire par_done_reg190_in;
  wire par_done_reg190_write_en;
  wire par_done_reg190_clk;
  wire par_done_reg190_out;
  wire par_done_reg190_done;
  wire par_done_reg191_in;
  wire par_done_reg191_write_en;
  wire par_done_reg191_clk;
  wire par_done_reg191_out;
  wire par_done_reg191_done;
  wire par_done_reg192_in;
  wire par_done_reg192_write_en;
  wire par_done_reg192_clk;
  wire par_done_reg192_out;
  wire par_done_reg192_done;
  wire par_done_reg193_in;
  wire par_done_reg193_write_en;
  wire par_done_reg193_clk;
  wire par_done_reg193_out;
  wire par_done_reg193_done;
  wire par_done_reg194_in;
  wire par_done_reg194_write_en;
  wire par_done_reg194_clk;
  wire par_done_reg194_out;
  wire par_done_reg194_done;
  wire par_done_reg195_in;
  wire par_done_reg195_write_en;
  wire par_done_reg195_clk;
  wire par_done_reg195_out;
  wire par_done_reg195_done;
  wire par_done_reg196_in;
  wire par_done_reg196_write_en;
  wire par_done_reg196_clk;
  wire par_done_reg196_out;
  wire par_done_reg196_done;
  wire par_done_reg197_in;
  wire par_done_reg197_write_en;
  wire par_done_reg197_clk;
  wire par_done_reg197_out;
  wire par_done_reg197_done;
  wire par_done_reg198_in;
  wire par_done_reg198_write_en;
  wire par_done_reg198_clk;
  wire par_done_reg198_out;
  wire par_done_reg198_done;
  wire par_done_reg199_in;
  wire par_done_reg199_write_en;
  wire par_done_reg199_clk;
  wire par_done_reg199_out;
  wire par_done_reg199_done;
  wire par_done_reg200_in;
  wire par_done_reg200_write_en;
  wire par_done_reg200_clk;
  wire par_done_reg200_out;
  wire par_done_reg200_done;
  wire par_done_reg201_in;
  wire par_done_reg201_write_en;
  wire par_done_reg201_clk;
  wire par_done_reg201_out;
  wire par_done_reg201_done;
  wire par_done_reg202_in;
  wire par_done_reg202_write_en;
  wire par_done_reg202_clk;
  wire par_done_reg202_out;
  wire par_done_reg202_done;
  wire par_done_reg203_in;
  wire par_done_reg203_write_en;
  wire par_done_reg203_clk;
  wire par_done_reg203_out;
  wire par_done_reg203_done;
  wire par_done_reg204_in;
  wire par_done_reg204_write_en;
  wire par_done_reg204_clk;
  wire par_done_reg204_out;
  wire par_done_reg204_done;
  wire par_done_reg205_in;
  wire par_done_reg205_write_en;
  wire par_done_reg205_clk;
  wire par_done_reg205_out;
  wire par_done_reg205_done;
  wire par_done_reg206_in;
  wire par_done_reg206_write_en;
  wire par_done_reg206_clk;
  wire par_done_reg206_out;
  wire par_done_reg206_done;
  wire par_done_reg207_in;
  wire par_done_reg207_write_en;
  wire par_done_reg207_clk;
  wire par_done_reg207_out;
  wire par_done_reg207_done;
  wire par_done_reg208_in;
  wire par_done_reg208_write_en;
  wire par_done_reg208_clk;
  wire par_done_reg208_out;
  wire par_done_reg208_done;
  wire par_done_reg209_in;
  wire par_done_reg209_write_en;
  wire par_done_reg209_clk;
  wire par_done_reg209_out;
  wire par_done_reg209_done;
  wire par_done_reg210_in;
  wire par_done_reg210_write_en;
  wire par_done_reg210_clk;
  wire par_done_reg210_out;
  wire par_done_reg210_done;
  wire par_done_reg211_in;
  wire par_done_reg211_write_en;
  wire par_done_reg211_clk;
  wire par_done_reg211_out;
  wire par_done_reg211_done;
  wire par_done_reg212_in;
  wire par_done_reg212_write_en;
  wire par_done_reg212_clk;
  wire par_done_reg212_out;
  wire par_done_reg212_done;
  wire par_reset14_in;
  wire par_reset14_write_en;
  wire par_reset14_clk;
  wire par_reset14_out;
  wire par_reset14_done;
  wire par_done_reg213_in;
  wire par_done_reg213_write_en;
  wire par_done_reg213_clk;
  wire par_done_reg213_out;
  wire par_done_reg213_done;
  wire par_done_reg214_in;
  wire par_done_reg214_write_en;
  wire par_done_reg214_clk;
  wire par_done_reg214_out;
  wire par_done_reg214_done;
  wire par_done_reg215_in;
  wire par_done_reg215_write_en;
  wire par_done_reg215_clk;
  wire par_done_reg215_out;
  wire par_done_reg215_done;
  wire par_done_reg216_in;
  wire par_done_reg216_write_en;
  wire par_done_reg216_clk;
  wire par_done_reg216_out;
  wire par_done_reg216_done;
  wire par_done_reg217_in;
  wire par_done_reg217_write_en;
  wire par_done_reg217_clk;
  wire par_done_reg217_out;
  wire par_done_reg217_done;
  wire par_done_reg218_in;
  wire par_done_reg218_write_en;
  wire par_done_reg218_clk;
  wire par_done_reg218_out;
  wire par_done_reg218_done;
  wire par_done_reg219_in;
  wire par_done_reg219_write_en;
  wire par_done_reg219_clk;
  wire par_done_reg219_out;
  wire par_done_reg219_done;
  wire par_done_reg220_in;
  wire par_done_reg220_write_en;
  wire par_done_reg220_clk;
  wire par_done_reg220_out;
  wire par_done_reg220_done;
  wire par_done_reg221_in;
  wire par_done_reg221_write_en;
  wire par_done_reg221_clk;
  wire par_done_reg221_out;
  wire par_done_reg221_done;
  wire par_done_reg222_in;
  wire par_done_reg222_write_en;
  wire par_done_reg222_clk;
  wire par_done_reg222_out;
  wire par_done_reg222_done;
  wire par_done_reg223_in;
  wire par_done_reg223_write_en;
  wire par_done_reg223_clk;
  wire par_done_reg223_out;
  wire par_done_reg223_done;
  wire par_done_reg224_in;
  wire par_done_reg224_write_en;
  wire par_done_reg224_clk;
  wire par_done_reg224_out;
  wire par_done_reg224_done;
  wire par_done_reg225_in;
  wire par_done_reg225_write_en;
  wire par_done_reg225_clk;
  wire par_done_reg225_out;
  wire par_done_reg225_done;
  wire par_done_reg226_in;
  wire par_done_reg226_write_en;
  wire par_done_reg226_clk;
  wire par_done_reg226_out;
  wire par_done_reg226_done;
  wire par_done_reg227_in;
  wire par_done_reg227_write_en;
  wire par_done_reg227_clk;
  wire par_done_reg227_out;
  wire par_done_reg227_done;
  wire par_done_reg228_in;
  wire par_done_reg228_write_en;
  wire par_done_reg228_clk;
  wire par_done_reg228_out;
  wire par_done_reg228_done;
  wire par_done_reg229_in;
  wire par_done_reg229_write_en;
  wire par_done_reg229_clk;
  wire par_done_reg229_out;
  wire par_done_reg229_done;
  wire par_done_reg230_in;
  wire par_done_reg230_write_en;
  wire par_done_reg230_clk;
  wire par_done_reg230_out;
  wire par_done_reg230_done;
  wire par_done_reg231_in;
  wire par_done_reg231_write_en;
  wire par_done_reg231_clk;
  wire par_done_reg231_out;
  wire par_done_reg231_done;
  wire par_done_reg232_in;
  wire par_done_reg232_write_en;
  wire par_done_reg232_clk;
  wire par_done_reg232_out;
  wire par_done_reg232_done;
  wire par_done_reg233_in;
  wire par_done_reg233_write_en;
  wire par_done_reg233_clk;
  wire par_done_reg233_out;
  wire par_done_reg233_done;
  wire par_done_reg234_in;
  wire par_done_reg234_write_en;
  wire par_done_reg234_clk;
  wire par_done_reg234_out;
  wire par_done_reg234_done;
  wire par_done_reg235_in;
  wire par_done_reg235_write_en;
  wire par_done_reg235_clk;
  wire par_done_reg235_out;
  wire par_done_reg235_done;
  wire par_done_reg236_in;
  wire par_done_reg236_write_en;
  wire par_done_reg236_clk;
  wire par_done_reg236_out;
  wire par_done_reg236_done;
  wire par_done_reg237_in;
  wire par_done_reg237_write_en;
  wire par_done_reg237_clk;
  wire par_done_reg237_out;
  wire par_done_reg237_done;
  wire par_done_reg238_in;
  wire par_done_reg238_write_en;
  wire par_done_reg238_clk;
  wire par_done_reg238_out;
  wire par_done_reg238_done;
  wire par_done_reg239_in;
  wire par_done_reg239_write_en;
  wire par_done_reg239_clk;
  wire par_done_reg239_out;
  wire par_done_reg239_done;
  wire par_done_reg240_in;
  wire par_done_reg240_write_en;
  wire par_done_reg240_clk;
  wire par_done_reg240_out;
  wire par_done_reg240_done;
  wire par_done_reg241_in;
  wire par_done_reg241_write_en;
  wire par_done_reg241_clk;
  wire par_done_reg241_out;
  wire par_done_reg241_done;
  wire par_done_reg242_in;
  wire par_done_reg242_write_en;
  wire par_done_reg242_clk;
  wire par_done_reg242_out;
  wire par_done_reg242_done;
  wire par_done_reg243_in;
  wire par_done_reg243_write_en;
  wire par_done_reg243_clk;
  wire par_done_reg243_out;
  wire par_done_reg243_done;
  wire par_done_reg244_in;
  wire par_done_reg244_write_en;
  wire par_done_reg244_clk;
  wire par_done_reg244_out;
  wire par_done_reg244_done;
  wire par_done_reg245_in;
  wire par_done_reg245_write_en;
  wire par_done_reg245_clk;
  wire par_done_reg245_out;
  wire par_done_reg245_done;
  wire par_done_reg246_in;
  wire par_done_reg246_write_en;
  wire par_done_reg246_clk;
  wire par_done_reg246_out;
  wire par_done_reg246_done;
  wire par_done_reg247_in;
  wire par_done_reg247_write_en;
  wire par_done_reg247_clk;
  wire par_done_reg247_out;
  wire par_done_reg247_done;
  wire par_done_reg248_in;
  wire par_done_reg248_write_en;
  wire par_done_reg248_clk;
  wire par_done_reg248_out;
  wire par_done_reg248_done;
  wire par_done_reg249_in;
  wire par_done_reg249_write_en;
  wire par_done_reg249_clk;
  wire par_done_reg249_out;
  wire par_done_reg249_done;
  wire par_done_reg250_in;
  wire par_done_reg250_write_en;
  wire par_done_reg250_clk;
  wire par_done_reg250_out;
  wire par_done_reg250_done;
  wire par_reset15_in;
  wire par_reset15_write_en;
  wire par_reset15_clk;
  wire par_reset15_out;
  wire par_reset15_done;
  wire par_done_reg251_in;
  wire par_done_reg251_write_en;
  wire par_done_reg251_clk;
  wire par_done_reg251_out;
  wire par_done_reg251_done;
  wire par_done_reg252_in;
  wire par_done_reg252_write_en;
  wire par_done_reg252_clk;
  wire par_done_reg252_out;
  wire par_done_reg252_done;
  wire par_done_reg253_in;
  wire par_done_reg253_write_en;
  wire par_done_reg253_clk;
  wire par_done_reg253_out;
  wire par_done_reg253_done;
  wire par_done_reg254_in;
  wire par_done_reg254_write_en;
  wire par_done_reg254_clk;
  wire par_done_reg254_out;
  wire par_done_reg254_done;
  wire par_done_reg255_in;
  wire par_done_reg255_write_en;
  wire par_done_reg255_clk;
  wire par_done_reg255_out;
  wire par_done_reg255_done;
  wire par_done_reg256_in;
  wire par_done_reg256_write_en;
  wire par_done_reg256_clk;
  wire par_done_reg256_out;
  wire par_done_reg256_done;
  wire par_done_reg257_in;
  wire par_done_reg257_write_en;
  wire par_done_reg257_clk;
  wire par_done_reg257_out;
  wire par_done_reg257_done;
  wire par_done_reg258_in;
  wire par_done_reg258_write_en;
  wire par_done_reg258_clk;
  wire par_done_reg258_out;
  wire par_done_reg258_done;
  wire par_done_reg259_in;
  wire par_done_reg259_write_en;
  wire par_done_reg259_clk;
  wire par_done_reg259_out;
  wire par_done_reg259_done;
  wire par_done_reg260_in;
  wire par_done_reg260_write_en;
  wire par_done_reg260_clk;
  wire par_done_reg260_out;
  wire par_done_reg260_done;
  wire par_done_reg261_in;
  wire par_done_reg261_write_en;
  wire par_done_reg261_clk;
  wire par_done_reg261_out;
  wire par_done_reg261_done;
  wire par_done_reg262_in;
  wire par_done_reg262_write_en;
  wire par_done_reg262_clk;
  wire par_done_reg262_out;
  wire par_done_reg262_done;
  wire par_done_reg263_in;
  wire par_done_reg263_write_en;
  wire par_done_reg263_clk;
  wire par_done_reg263_out;
  wire par_done_reg263_done;
  wire par_done_reg264_in;
  wire par_done_reg264_write_en;
  wire par_done_reg264_clk;
  wire par_done_reg264_out;
  wire par_done_reg264_done;
  wire par_done_reg265_in;
  wire par_done_reg265_write_en;
  wire par_done_reg265_clk;
  wire par_done_reg265_out;
  wire par_done_reg265_done;
  wire par_done_reg266_in;
  wire par_done_reg266_write_en;
  wire par_done_reg266_clk;
  wire par_done_reg266_out;
  wire par_done_reg266_done;
  wire par_done_reg267_in;
  wire par_done_reg267_write_en;
  wire par_done_reg267_clk;
  wire par_done_reg267_out;
  wire par_done_reg267_done;
  wire par_done_reg268_in;
  wire par_done_reg268_write_en;
  wire par_done_reg268_clk;
  wire par_done_reg268_out;
  wire par_done_reg268_done;
  wire par_done_reg269_in;
  wire par_done_reg269_write_en;
  wire par_done_reg269_clk;
  wire par_done_reg269_out;
  wire par_done_reg269_done;
  wire par_done_reg270_in;
  wire par_done_reg270_write_en;
  wire par_done_reg270_clk;
  wire par_done_reg270_out;
  wire par_done_reg270_done;
  wire par_done_reg271_in;
  wire par_done_reg271_write_en;
  wire par_done_reg271_clk;
  wire par_done_reg271_out;
  wire par_done_reg271_done;
  wire par_done_reg272_in;
  wire par_done_reg272_write_en;
  wire par_done_reg272_clk;
  wire par_done_reg272_out;
  wire par_done_reg272_done;
  wire par_done_reg273_in;
  wire par_done_reg273_write_en;
  wire par_done_reg273_clk;
  wire par_done_reg273_out;
  wire par_done_reg273_done;
  wire par_reset16_in;
  wire par_reset16_write_en;
  wire par_reset16_clk;
  wire par_reset16_out;
  wire par_reset16_done;
  wire par_done_reg274_in;
  wire par_done_reg274_write_en;
  wire par_done_reg274_clk;
  wire par_done_reg274_out;
  wire par_done_reg274_done;
  wire par_done_reg275_in;
  wire par_done_reg275_write_en;
  wire par_done_reg275_clk;
  wire par_done_reg275_out;
  wire par_done_reg275_done;
  wire par_done_reg276_in;
  wire par_done_reg276_write_en;
  wire par_done_reg276_clk;
  wire par_done_reg276_out;
  wire par_done_reg276_done;
  wire par_done_reg277_in;
  wire par_done_reg277_write_en;
  wire par_done_reg277_clk;
  wire par_done_reg277_out;
  wire par_done_reg277_done;
  wire par_done_reg278_in;
  wire par_done_reg278_write_en;
  wire par_done_reg278_clk;
  wire par_done_reg278_out;
  wire par_done_reg278_done;
  wire par_done_reg279_in;
  wire par_done_reg279_write_en;
  wire par_done_reg279_clk;
  wire par_done_reg279_out;
  wire par_done_reg279_done;
  wire par_done_reg280_in;
  wire par_done_reg280_write_en;
  wire par_done_reg280_clk;
  wire par_done_reg280_out;
  wire par_done_reg280_done;
  wire par_done_reg281_in;
  wire par_done_reg281_write_en;
  wire par_done_reg281_clk;
  wire par_done_reg281_out;
  wire par_done_reg281_done;
  wire par_done_reg282_in;
  wire par_done_reg282_write_en;
  wire par_done_reg282_clk;
  wire par_done_reg282_out;
  wire par_done_reg282_done;
  wire par_done_reg283_in;
  wire par_done_reg283_write_en;
  wire par_done_reg283_clk;
  wire par_done_reg283_out;
  wire par_done_reg283_done;
  wire par_done_reg284_in;
  wire par_done_reg284_write_en;
  wire par_done_reg284_clk;
  wire par_done_reg284_out;
  wire par_done_reg284_done;
  wire par_done_reg285_in;
  wire par_done_reg285_write_en;
  wire par_done_reg285_clk;
  wire par_done_reg285_out;
  wire par_done_reg285_done;
  wire par_done_reg286_in;
  wire par_done_reg286_write_en;
  wire par_done_reg286_clk;
  wire par_done_reg286_out;
  wire par_done_reg286_done;
  wire par_done_reg287_in;
  wire par_done_reg287_write_en;
  wire par_done_reg287_clk;
  wire par_done_reg287_out;
  wire par_done_reg287_done;
  wire par_done_reg288_in;
  wire par_done_reg288_write_en;
  wire par_done_reg288_clk;
  wire par_done_reg288_out;
  wire par_done_reg288_done;
  wire par_done_reg289_in;
  wire par_done_reg289_write_en;
  wire par_done_reg289_clk;
  wire par_done_reg289_out;
  wire par_done_reg289_done;
  wire par_done_reg290_in;
  wire par_done_reg290_write_en;
  wire par_done_reg290_clk;
  wire par_done_reg290_out;
  wire par_done_reg290_done;
  wire par_done_reg291_in;
  wire par_done_reg291_write_en;
  wire par_done_reg291_clk;
  wire par_done_reg291_out;
  wire par_done_reg291_done;
  wire par_done_reg292_in;
  wire par_done_reg292_write_en;
  wire par_done_reg292_clk;
  wire par_done_reg292_out;
  wire par_done_reg292_done;
  wire par_done_reg293_in;
  wire par_done_reg293_write_en;
  wire par_done_reg293_clk;
  wire par_done_reg293_out;
  wire par_done_reg293_done;
  wire par_done_reg294_in;
  wire par_done_reg294_write_en;
  wire par_done_reg294_clk;
  wire par_done_reg294_out;
  wire par_done_reg294_done;
  wire par_done_reg295_in;
  wire par_done_reg295_write_en;
  wire par_done_reg295_clk;
  wire par_done_reg295_out;
  wire par_done_reg295_done;
  wire par_done_reg296_in;
  wire par_done_reg296_write_en;
  wire par_done_reg296_clk;
  wire par_done_reg296_out;
  wire par_done_reg296_done;
  wire par_done_reg297_in;
  wire par_done_reg297_write_en;
  wire par_done_reg297_clk;
  wire par_done_reg297_out;
  wire par_done_reg297_done;
  wire par_done_reg298_in;
  wire par_done_reg298_write_en;
  wire par_done_reg298_clk;
  wire par_done_reg298_out;
  wire par_done_reg298_done;
  wire par_done_reg299_in;
  wire par_done_reg299_write_en;
  wire par_done_reg299_clk;
  wire par_done_reg299_out;
  wire par_done_reg299_done;
  wire par_done_reg300_in;
  wire par_done_reg300_write_en;
  wire par_done_reg300_clk;
  wire par_done_reg300_out;
  wire par_done_reg300_done;
  wire par_done_reg301_in;
  wire par_done_reg301_write_en;
  wire par_done_reg301_clk;
  wire par_done_reg301_out;
  wire par_done_reg301_done;
  wire par_done_reg302_in;
  wire par_done_reg302_write_en;
  wire par_done_reg302_clk;
  wire par_done_reg302_out;
  wire par_done_reg302_done;
  wire par_done_reg303_in;
  wire par_done_reg303_write_en;
  wire par_done_reg303_clk;
  wire par_done_reg303_out;
  wire par_done_reg303_done;
  wire par_done_reg304_in;
  wire par_done_reg304_write_en;
  wire par_done_reg304_clk;
  wire par_done_reg304_out;
  wire par_done_reg304_done;
  wire par_done_reg305_in;
  wire par_done_reg305_write_en;
  wire par_done_reg305_clk;
  wire par_done_reg305_out;
  wire par_done_reg305_done;
  wire par_done_reg306_in;
  wire par_done_reg306_write_en;
  wire par_done_reg306_clk;
  wire par_done_reg306_out;
  wire par_done_reg306_done;
  wire par_done_reg307_in;
  wire par_done_reg307_write_en;
  wire par_done_reg307_clk;
  wire par_done_reg307_out;
  wire par_done_reg307_done;
  wire par_done_reg308_in;
  wire par_done_reg308_write_en;
  wire par_done_reg308_clk;
  wire par_done_reg308_out;
  wire par_done_reg308_done;
  wire par_done_reg309_in;
  wire par_done_reg309_write_en;
  wire par_done_reg309_clk;
  wire par_done_reg309_out;
  wire par_done_reg309_done;
  wire par_reset17_in;
  wire par_reset17_write_en;
  wire par_reset17_clk;
  wire par_reset17_out;
  wire par_reset17_done;
  wire par_done_reg310_in;
  wire par_done_reg310_write_en;
  wire par_done_reg310_clk;
  wire par_done_reg310_out;
  wire par_done_reg310_done;
  wire par_done_reg311_in;
  wire par_done_reg311_write_en;
  wire par_done_reg311_clk;
  wire par_done_reg311_out;
  wire par_done_reg311_done;
  wire par_done_reg312_in;
  wire par_done_reg312_write_en;
  wire par_done_reg312_clk;
  wire par_done_reg312_out;
  wire par_done_reg312_done;
  wire par_done_reg313_in;
  wire par_done_reg313_write_en;
  wire par_done_reg313_clk;
  wire par_done_reg313_out;
  wire par_done_reg313_done;
  wire par_done_reg314_in;
  wire par_done_reg314_write_en;
  wire par_done_reg314_clk;
  wire par_done_reg314_out;
  wire par_done_reg314_done;
  wire par_done_reg315_in;
  wire par_done_reg315_write_en;
  wire par_done_reg315_clk;
  wire par_done_reg315_out;
  wire par_done_reg315_done;
  wire par_done_reg316_in;
  wire par_done_reg316_write_en;
  wire par_done_reg316_clk;
  wire par_done_reg316_out;
  wire par_done_reg316_done;
  wire par_done_reg317_in;
  wire par_done_reg317_write_en;
  wire par_done_reg317_clk;
  wire par_done_reg317_out;
  wire par_done_reg317_done;
  wire par_done_reg318_in;
  wire par_done_reg318_write_en;
  wire par_done_reg318_clk;
  wire par_done_reg318_out;
  wire par_done_reg318_done;
  wire par_done_reg319_in;
  wire par_done_reg319_write_en;
  wire par_done_reg319_clk;
  wire par_done_reg319_out;
  wire par_done_reg319_done;
  wire par_done_reg320_in;
  wire par_done_reg320_write_en;
  wire par_done_reg320_clk;
  wire par_done_reg320_out;
  wire par_done_reg320_done;
  wire par_done_reg321_in;
  wire par_done_reg321_write_en;
  wire par_done_reg321_clk;
  wire par_done_reg321_out;
  wire par_done_reg321_done;
  wire par_done_reg322_in;
  wire par_done_reg322_write_en;
  wire par_done_reg322_clk;
  wire par_done_reg322_out;
  wire par_done_reg322_done;
  wire par_done_reg323_in;
  wire par_done_reg323_write_en;
  wire par_done_reg323_clk;
  wire par_done_reg323_out;
  wire par_done_reg323_done;
  wire par_done_reg324_in;
  wire par_done_reg324_write_en;
  wire par_done_reg324_clk;
  wire par_done_reg324_out;
  wire par_done_reg324_done;
  wire par_done_reg325_in;
  wire par_done_reg325_write_en;
  wire par_done_reg325_clk;
  wire par_done_reg325_out;
  wire par_done_reg325_done;
  wire par_done_reg326_in;
  wire par_done_reg326_write_en;
  wire par_done_reg326_clk;
  wire par_done_reg326_out;
  wire par_done_reg326_done;
  wire par_done_reg327_in;
  wire par_done_reg327_write_en;
  wire par_done_reg327_clk;
  wire par_done_reg327_out;
  wire par_done_reg327_done;
  wire par_done_reg328_in;
  wire par_done_reg328_write_en;
  wire par_done_reg328_clk;
  wire par_done_reg328_out;
  wire par_done_reg328_done;
  wire par_done_reg329_in;
  wire par_done_reg329_write_en;
  wire par_done_reg329_clk;
  wire par_done_reg329_out;
  wire par_done_reg329_done;
  wire par_reset18_in;
  wire par_reset18_write_en;
  wire par_reset18_clk;
  wire par_reset18_out;
  wire par_reset18_done;
  wire par_done_reg330_in;
  wire par_done_reg330_write_en;
  wire par_done_reg330_clk;
  wire par_done_reg330_out;
  wire par_done_reg330_done;
  wire par_done_reg331_in;
  wire par_done_reg331_write_en;
  wire par_done_reg331_clk;
  wire par_done_reg331_out;
  wire par_done_reg331_done;
  wire par_done_reg332_in;
  wire par_done_reg332_write_en;
  wire par_done_reg332_clk;
  wire par_done_reg332_out;
  wire par_done_reg332_done;
  wire par_done_reg333_in;
  wire par_done_reg333_write_en;
  wire par_done_reg333_clk;
  wire par_done_reg333_out;
  wire par_done_reg333_done;
  wire par_done_reg334_in;
  wire par_done_reg334_write_en;
  wire par_done_reg334_clk;
  wire par_done_reg334_out;
  wire par_done_reg334_done;
  wire par_done_reg335_in;
  wire par_done_reg335_write_en;
  wire par_done_reg335_clk;
  wire par_done_reg335_out;
  wire par_done_reg335_done;
  wire par_done_reg336_in;
  wire par_done_reg336_write_en;
  wire par_done_reg336_clk;
  wire par_done_reg336_out;
  wire par_done_reg336_done;
  wire par_done_reg337_in;
  wire par_done_reg337_write_en;
  wire par_done_reg337_clk;
  wire par_done_reg337_out;
  wire par_done_reg337_done;
  wire par_done_reg338_in;
  wire par_done_reg338_write_en;
  wire par_done_reg338_clk;
  wire par_done_reg338_out;
  wire par_done_reg338_done;
  wire par_done_reg339_in;
  wire par_done_reg339_write_en;
  wire par_done_reg339_clk;
  wire par_done_reg339_out;
  wire par_done_reg339_done;
  wire par_done_reg340_in;
  wire par_done_reg340_write_en;
  wire par_done_reg340_clk;
  wire par_done_reg340_out;
  wire par_done_reg340_done;
  wire par_done_reg341_in;
  wire par_done_reg341_write_en;
  wire par_done_reg341_clk;
  wire par_done_reg341_out;
  wire par_done_reg341_done;
  wire par_done_reg342_in;
  wire par_done_reg342_write_en;
  wire par_done_reg342_clk;
  wire par_done_reg342_out;
  wire par_done_reg342_done;
  wire par_done_reg343_in;
  wire par_done_reg343_write_en;
  wire par_done_reg343_clk;
  wire par_done_reg343_out;
  wire par_done_reg343_done;
  wire par_done_reg344_in;
  wire par_done_reg344_write_en;
  wire par_done_reg344_clk;
  wire par_done_reg344_out;
  wire par_done_reg344_done;
  wire par_done_reg345_in;
  wire par_done_reg345_write_en;
  wire par_done_reg345_clk;
  wire par_done_reg345_out;
  wire par_done_reg345_done;
  wire par_done_reg346_in;
  wire par_done_reg346_write_en;
  wire par_done_reg346_clk;
  wire par_done_reg346_out;
  wire par_done_reg346_done;
  wire par_done_reg347_in;
  wire par_done_reg347_write_en;
  wire par_done_reg347_clk;
  wire par_done_reg347_out;
  wire par_done_reg347_done;
  wire par_done_reg348_in;
  wire par_done_reg348_write_en;
  wire par_done_reg348_clk;
  wire par_done_reg348_out;
  wire par_done_reg348_done;
  wire par_done_reg349_in;
  wire par_done_reg349_write_en;
  wire par_done_reg349_clk;
  wire par_done_reg349_out;
  wire par_done_reg349_done;
  wire par_done_reg350_in;
  wire par_done_reg350_write_en;
  wire par_done_reg350_clk;
  wire par_done_reg350_out;
  wire par_done_reg350_done;
  wire par_done_reg351_in;
  wire par_done_reg351_write_en;
  wire par_done_reg351_clk;
  wire par_done_reg351_out;
  wire par_done_reg351_done;
  wire par_done_reg352_in;
  wire par_done_reg352_write_en;
  wire par_done_reg352_clk;
  wire par_done_reg352_out;
  wire par_done_reg352_done;
  wire par_done_reg353_in;
  wire par_done_reg353_write_en;
  wire par_done_reg353_clk;
  wire par_done_reg353_out;
  wire par_done_reg353_done;
  wire par_done_reg354_in;
  wire par_done_reg354_write_en;
  wire par_done_reg354_clk;
  wire par_done_reg354_out;
  wire par_done_reg354_done;
  wire par_done_reg355_in;
  wire par_done_reg355_write_en;
  wire par_done_reg355_clk;
  wire par_done_reg355_out;
  wire par_done_reg355_done;
  wire par_done_reg356_in;
  wire par_done_reg356_write_en;
  wire par_done_reg356_clk;
  wire par_done_reg356_out;
  wire par_done_reg356_done;
  wire par_done_reg357_in;
  wire par_done_reg357_write_en;
  wire par_done_reg357_clk;
  wire par_done_reg357_out;
  wire par_done_reg357_done;
  wire par_done_reg358_in;
  wire par_done_reg358_write_en;
  wire par_done_reg358_clk;
  wire par_done_reg358_out;
  wire par_done_reg358_done;
  wire par_done_reg359_in;
  wire par_done_reg359_write_en;
  wire par_done_reg359_clk;
  wire par_done_reg359_out;
  wire par_done_reg359_done;
  wire par_reset19_in;
  wire par_reset19_write_en;
  wire par_reset19_clk;
  wire par_reset19_out;
  wire par_reset19_done;
  wire par_done_reg360_in;
  wire par_done_reg360_write_en;
  wire par_done_reg360_clk;
  wire par_done_reg360_out;
  wire par_done_reg360_done;
  wire par_done_reg361_in;
  wire par_done_reg361_write_en;
  wire par_done_reg361_clk;
  wire par_done_reg361_out;
  wire par_done_reg361_done;
  wire par_done_reg362_in;
  wire par_done_reg362_write_en;
  wire par_done_reg362_clk;
  wire par_done_reg362_out;
  wire par_done_reg362_done;
  wire par_done_reg363_in;
  wire par_done_reg363_write_en;
  wire par_done_reg363_clk;
  wire par_done_reg363_out;
  wire par_done_reg363_done;
  wire par_done_reg364_in;
  wire par_done_reg364_write_en;
  wire par_done_reg364_clk;
  wire par_done_reg364_out;
  wire par_done_reg364_done;
  wire par_done_reg365_in;
  wire par_done_reg365_write_en;
  wire par_done_reg365_clk;
  wire par_done_reg365_out;
  wire par_done_reg365_done;
  wire par_done_reg366_in;
  wire par_done_reg366_write_en;
  wire par_done_reg366_clk;
  wire par_done_reg366_out;
  wire par_done_reg366_done;
  wire par_done_reg367_in;
  wire par_done_reg367_write_en;
  wire par_done_reg367_clk;
  wire par_done_reg367_out;
  wire par_done_reg367_done;
  wire par_done_reg368_in;
  wire par_done_reg368_write_en;
  wire par_done_reg368_clk;
  wire par_done_reg368_out;
  wire par_done_reg368_done;
  wire par_done_reg369_in;
  wire par_done_reg369_write_en;
  wire par_done_reg369_clk;
  wire par_done_reg369_out;
  wire par_done_reg369_done;
  wire par_done_reg370_in;
  wire par_done_reg370_write_en;
  wire par_done_reg370_clk;
  wire par_done_reg370_out;
  wire par_done_reg370_done;
  wire par_done_reg371_in;
  wire par_done_reg371_write_en;
  wire par_done_reg371_clk;
  wire par_done_reg371_out;
  wire par_done_reg371_done;
  wire par_done_reg372_in;
  wire par_done_reg372_write_en;
  wire par_done_reg372_clk;
  wire par_done_reg372_out;
  wire par_done_reg372_done;
  wire par_done_reg373_in;
  wire par_done_reg373_write_en;
  wire par_done_reg373_clk;
  wire par_done_reg373_out;
  wire par_done_reg373_done;
  wire par_done_reg374_in;
  wire par_done_reg374_write_en;
  wire par_done_reg374_clk;
  wire par_done_reg374_out;
  wire par_done_reg374_done;
  wire par_reset20_in;
  wire par_reset20_write_en;
  wire par_reset20_clk;
  wire par_reset20_out;
  wire par_reset20_done;
  wire par_done_reg375_in;
  wire par_done_reg375_write_en;
  wire par_done_reg375_clk;
  wire par_done_reg375_out;
  wire par_done_reg375_done;
  wire par_done_reg376_in;
  wire par_done_reg376_write_en;
  wire par_done_reg376_clk;
  wire par_done_reg376_out;
  wire par_done_reg376_done;
  wire par_done_reg377_in;
  wire par_done_reg377_write_en;
  wire par_done_reg377_clk;
  wire par_done_reg377_out;
  wire par_done_reg377_done;
  wire par_done_reg378_in;
  wire par_done_reg378_write_en;
  wire par_done_reg378_clk;
  wire par_done_reg378_out;
  wire par_done_reg378_done;
  wire par_done_reg379_in;
  wire par_done_reg379_write_en;
  wire par_done_reg379_clk;
  wire par_done_reg379_out;
  wire par_done_reg379_done;
  wire par_done_reg380_in;
  wire par_done_reg380_write_en;
  wire par_done_reg380_clk;
  wire par_done_reg380_out;
  wire par_done_reg380_done;
  wire par_done_reg381_in;
  wire par_done_reg381_write_en;
  wire par_done_reg381_clk;
  wire par_done_reg381_out;
  wire par_done_reg381_done;
  wire par_done_reg382_in;
  wire par_done_reg382_write_en;
  wire par_done_reg382_clk;
  wire par_done_reg382_out;
  wire par_done_reg382_done;
  wire par_done_reg383_in;
  wire par_done_reg383_write_en;
  wire par_done_reg383_clk;
  wire par_done_reg383_out;
  wire par_done_reg383_done;
  wire par_done_reg384_in;
  wire par_done_reg384_write_en;
  wire par_done_reg384_clk;
  wire par_done_reg384_out;
  wire par_done_reg384_done;
  wire par_done_reg385_in;
  wire par_done_reg385_write_en;
  wire par_done_reg385_clk;
  wire par_done_reg385_out;
  wire par_done_reg385_done;
  wire par_done_reg386_in;
  wire par_done_reg386_write_en;
  wire par_done_reg386_clk;
  wire par_done_reg386_out;
  wire par_done_reg386_done;
  wire par_done_reg387_in;
  wire par_done_reg387_write_en;
  wire par_done_reg387_clk;
  wire par_done_reg387_out;
  wire par_done_reg387_done;
  wire par_done_reg388_in;
  wire par_done_reg388_write_en;
  wire par_done_reg388_clk;
  wire par_done_reg388_out;
  wire par_done_reg388_done;
  wire par_done_reg389_in;
  wire par_done_reg389_write_en;
  wire par_done_reg389_clk;
  wire par_done_reg389_out;
  wire par_done_reg389_done;
  wire par_done_reg390_in;
  wire par_done_reg390_write_en;
  wire par_done_reg390_clk;
  wire par_done_reg390_out;
  wire par_done_reg390_done;
  wire par_done_reg391_in;
  wire par_done_reg391_write_en;
  wire par_done_reg391_clk;
  wire par_done_reg391_out;
  wire par_done_reg391_done;
  wire par_done_reg392_in;
  wire par_done_reg392_write_en;
  wire par_done_reg392_clk;
  wire par_done_reg392_out;
  wire par_done_reg392_done;
  wire par_done_reg393_in;
  wire par_done_reg393_write_en;
  wire par_done_reg393_clk;
  wire par_done_reg393_out;
  wire par_done_reg393_done;
  wire par_done_reg394_in;
  wire par_done_reg394_write_en;
  wire par_done_reg394_clk;
  wire par_done_reg394_out;
  wire par_done_reg394_done;
  wire par_reset21_in;
  wire par_reset21_write_en;
  wire par_reset21_clk;
  wire par_reset21_out;
  wire par_reset21_done;
  wire par_done_reg395_in;
  wire par_done_reg395_write_en;
  wire par_done_reg395_clk;
  wire par_done_reg395_out;
  wire par_done_reg395_done;
  wire par_done_reg396_in;
  wire par_done_reg396_write_en;
  wire par_done_reg396_clk;
  wire par_done_reg396_out;
  wire par_done_reg396_done;
  wire par_done_reg397_in;
  wire par_done_reg397_write_en;
  wire par_done_reg397_clk;
  wire par_done_reg397_out;
  wire par_done_reg397_done;
  wire par_done_reg398_in;
  wire par_done_reg398_write_en;
  wire par_done_reg398_clk;
  wire par_done_reg398_out;
  wire par_done_reg398_done;
  wire par_done_reg399_in;
  wire par_done_reg399_write_en;
  wire par_done_reg399_clk;
  wire par_done_reg399_out;
  wire par_done_reg399_done;
  wire par_done_reg400_in;
  wire par_done_reg400_write_en;
  wire par_done_reg400_clk;
  wire par_done_reg400_out;
  wire par_done_reg400_done;
  wire par_done_reg401_in;
  wire par_done_reg401_write_en;
  wire par_done_reg401_clk;
  wire par_done_reg401_out;
  wire par_done_reg401_done;
  wire par_done_reg402_in;
  wire par_done_reg402_write_en;
  wire par_done_reg402_clk;
  wire par_done_reg402_out;
  wire par_done_reg402_done;
  wire par_done_reg403_in;
  wire par_done_reg403_write_en;
  wire par_done_reg403_clk;
  wire par_done_reg403_out;
  wire par_done_reg403_done;
  wire par_done_reg404_in;
  wire par_done_reg404_write_en;
  wire par_done_reg404_clk;
  wire par_done_reg404_out;
  wire par_done_reg404_done;
  wire par_reset22_in;
  wire par_reset22_write_en;
  wire par_reset22_clk;
  wire par_reset22_out;
  wire par_reset22_done;
  wire par_done_reg405_in;
  wire par_done_reg405_write_en;
  wire par_done_reg405_clk;
  wire par_done_reg405_out;
  wire par_done_reg405_done;
  wire par_done_reg406_in;
  wire par_done_reg406_write_en;
  wire par_done_reg406_clk;
  wire par_done_reg406_out;
  wire par_done_reg406_done;
  wire par_done_reg407_in;
  wire par_done_reg407_write_en;
  wire par_done_reg407_clk;
  wire par_done_reg407_out;
  wire par_done_reg407_done;
  wire par_done_reg408_in;
  wire par_done_reg408_write_en;
  wire par_done_reg408_clk;
  wire par_done_reg408_out;
  wire par_done_reg408_done;
  wire par_done_reg409_in;
  wire par_done_reg409_write_en;
  wire par_done_reg409_clk;
  wire par_done_reg409_out;
  wire par_done_reg409_done;
  wire par_done_reg410_in;
  wire par_done_reg410_write_en;
  wire par_done_reg410_clk;
  wire par_done_reg410_out;
  wire par_done_reg410_done;
  wire par_done_reg411_in;
  wire par_done_reg411_write_en;
  wire par_done_reg411_clk;
  wire par_done_reg411_out;
  wire par_done_reg411_done;
  wire par_done_reg412_in;
  wire par_done_reg412_write_en;
  wire par_done_reg412_clk;
  wire par_done_reg412_out;
  wire par_done_reg412_done;
  wire par_done_reg413_in;
  wire par_done_reg413_write_en;
  wire par_done_reg413_clk;
  wire par_done_reg413_out;
  wire par_done_reg413_done;
  wire par_done_reg414_in;
  wire par_done_reg414_write_en;
  wire par_done_reg414_clk;
  wire par_done_reg414_out;
  wire par_done_reg414_done;
  wire par_done_reg415_in;
  wire par_done_reg415_write_en;
  wire par_done_reg415_clk;
  wire par_done_reg415_out;
  wire par_done_reg415_done;
  wire par_done_reg416_in;
  wire par_done_reg416_write_en;
  wire par_done_reg416_clk;
  wire par_done_reg416_out;
  wire par_done_reg416_done;
  wire par_reset23_in;
  wire par_reset23_write_en;
  wire par_reset23_clk;
  wire par_reset23_out;
  wire par_reset23_done;
  wire par_done_reg417_in;
  wire par_done_reg417_write_en;
  wire par_done_reg417_clk;
  wire par_done_reg417_out;
  wire par_done_reg417_done;
  wire par_done_reg418_in;
  wire par_done_reg418_write_en;
  wire par_done_reg418_clk;
  wire par_done_reg418_out;
  wire par_done_reg418_done;
  wire par_done_reg419_in;
  wire par_done_reg419_write_en;
  wire par_done_reg419_clk;
  wire par_done_reg419_out;
  wire par_done_reg419_done;
  wire par_done_reg420_in;
  wire par_done_reg420_write_en;
  wire par_done_reg420_clk;
  wire par_done_reg420_out;
  wire par_done_reg420_done;
  wire par_done_reg421_in;
  wire par_done_reg421_write_en;
  wire par_done_reg421_clk;
  wire par_done_reg421_out;
  wire par_done_reg421_done;
  wire par_done_reg422_in;
  wire par_done_reg422_write_en;
  wire par_done_reg422_clk;
  wire par_done_reg422_out;
  wire par_done_reg422_done;
  wire par_reset24_in;
  wire par_reset24_write_en;
  wire par_reset24_clk;
  wire par_reset24_out;
  wire par_reset24_done;
  wire par_done_reg423_in;
  wire par_done_reg423_write_en;
  wire par_done_reg423_clk;
  wire par_done_reg423_out;
  wire par_done_reg423_done;
  wire par_done_reg424_in;
  wire par_done_reg424_write_en;
  wire par_done_reg424_clk;
  wire par_done_reg424_out;
  wire par_done_reg424_done;
  wire par_done_reg425_in;
  wire par_done_reg425_write_en;
  wire par_done_reg425_clk;
  wire par_done_reg425_out;
  wire par_done_reg425_done;
  wire par_done_reg426_in;
  wire par_done_reg426_write_en;
  wire par_done_reg426_clk;
  wire par_done_reg426_out;
  wire par_done_reg426_done;
  wire par_done_reg427_in;
  wire par_done_reg427_write_en;
  wire par_done_reg427_clk;
  wire par_done_reg427_out;
  wire par_done_reg427_done;
  wire par_done_reg428_in;
  wire par_done_reg428_write_en;
  wire par_done_reg428_clk;
  wire par_done_reg428_out;
  wire par_done_reg428_done;
  wire par_reset25_in;
  wire par_reset25_write_en;
  wire par_reset25_clk;
  wire par_reset25_out;
  wire par_reset25_done;
  wire par_done_reg429_in;
  wire par_done_reg429_write_en;
  wire par_done_reg429_clk;
  wire par_done_reg429_out;
  wire par_done_reg429_done;
  wire par_done_reg430_in;
  wire par_done_reg430_write_en;
  wire par_done_reg430_clk;
  wire par_done_reg430_out;
  wire par_done_reg430_done;
  wire par_done_reg431_in;
  wire par_done_reg431_write_en;
  wire par_done_reg431_clk;
  wire par_done_reg431_out;
  wire par_done_reg431_done;
  wire par_reset26_in;
  wire par_reset26_write_en;
  wire par_reset26_clk;
  wire par_reset26_out;
  wire par_reset26_done;
  wire par_done_reg432_in;
  wire par_done_reg432_write_en;
  wire par_done_reg432_clk;
  wire par_done_reg432_out;
  wire par_done_reg432_done;
  wire par_done_reg433_in;
  wire par_done_reg433_write_en;
  wire par_done_reg433_clk;
  wire par_done_reg433_out;
  wire par_done_reg433_done;
  wire par_reset27_in;
  wire par_reset27_write_en;
  wire par_reset27_clk;
  wire par_reset27_out;
  wire par_reset27_done;
  wire par_done_reg434_in;
  wire par_done_reg434_write_en;
  wire par_done_reg434_clk;
  wire par_done_reg434_out;
  wire par_done_reg434_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_reg #(32) left_44_read (
      .in(left_44_read_in),
      .write_en(left_44_read_write_en),
      .clk(clk),
      .out(left_44_read_out),
      .done(left_44_read_done)
  );
  
  std_reg #(32) top_44_read (
      .in(top_44_read_in),
      .write_en(top_44_read_write_en),
      .clk(clk),
      .out(top_44_read_out),
      .done(top_44_read_done)
  );
  
  mac_pe #() pe_44 (
      .top(pe_44_top),
      .left(pe_44_left),
      .go(pe_44_go),
      .clk(clk),
      .down(pe_44_down),
      .right(pe_44_right),
      .out(pe_44_out),
      .done(pe_44_done)
  );
  
  std_reg #(32) right_43_write (
      .in(right_43_write_in),
      .write_en(right_43_write_write_en),
      .clk(clk),
      .out(right_43_write_out),
      .done(right_43_write_done)
  );
  
  std_reg #(32) left_43_read (
      .in(left_43_read_in),
      .write_en(left_43_read_write_en),
      .clk(clk),
      .out(left_43_read_out),
      .done(left_43_read_done)
  );
  
  std_reg #(32) top_43_read (
      .in(top_43_read_in),
      .write_en(top_43_read_write_en),
      .clk(clk),
      .out(top_43_read_out),
      .done(top_43_read_done)
  );
  
  mac_pe #() pe_43 (
      .top(pe_43_top),
      .left(pe_43_left),
      .go(pe_43_go),
      .clk(clk),
      .down(pe_43_down),
      .right(pe_43_right),
      .out(pe_43_out),
      .done(pe_43_done)
  );
  
  std_reg #(32) right_42_write (
      .in(right_42_write_in),
      .write_en(right_42_write_write_en),
      .clk(clk),
      .out(right_42_write_out),
      .done(right_42_write_done)
  );
  
  std_reg #(32) left_42_read (
      .in(left_42_read_in),
      .write_en(left_42_read_write_en),
      .clk(clk),
      .out(left_42_read_out),
      .done(left_42_read_done)
  );
  
  std_reg #(32) top_42_read (
      .in(top_42_read_in),
      .write_en(top_42_read_write_en),
      .clk(clk),
      .out(top_42_read_out),
      .done(top_42_read_done)
  );
  
  mac_pe #() pe_42 (
      .top(pe_42_top),
      .left(pe_42_left),
      .go(pe_42_go),
      .clk(clk),
      .down(pe_42_down),
      .right(pe_42_right),
      .out(pe_42_out),
      .done(pe_42_done)
  );
  
  std_reg #(32) right_41_write (
      .in(right_41_write_in),
      .write_en(right_41_write_write_en),
      .clk(clk),
      .out(right_41_write_out),
      .done(right_41_write_done)
  );
  
  std_reg #(32) left_41_read (
      .in(left_41_read_in),
      .write_en(left_41_read_write_en),
      .clk(clk),
      .out(left_41_read_out),
      .done(left_41_read_done)
  );
  
  std_reg #(32) top_41_read (
      .in(top_41_read_in),
      .write_en(top_41_read_write_en),
      .clk(clk),
      .out(top_41_read_out),
      .done(top_41_read_done)
  );
  
  mac_pe #() pe_41 (
      .top(pe_41_top),
      .left(pe_41_left),
      .go(pe_41_go),
      .clk(clk),
      .down(pe_41_down),
      .right(pe_41_right),
      .out(pe_41_out),
      .done(pe_41_done)
  );
  
  std_reg #(32) right_40_write (
      .in(right_40_write_in),
      .write_en(right_40_write_write_en),
      .clk(clk),
      .out(right_40_write_out),
      .done(right_40_write_done)
  );
  
  std_reg #(32) left_40_read (
      .in(left_40_read_in),
      .write_en(left_40_read_write_en),
      .clk(clk),
      .out(left_40_read_out),
      .done(left_40_read_done)
  );
  
  std_reg #(32) top_40_read (
      .in(top_40_read_in),
      .write_en(top_40_read_write_en),
      .clk(clk),
      .out(top_40_read_out),
      .done(top_40_read_done)
  );
  
  mac_pe #() pe_40 (
      .top(pe_40_top),
      .left(pe_40_left),
      .go(pe_40_go),
      .clk(clk),
      .down(pe_40_down),
      .right(pe_40_right),
      .out(pe_40_out),
      .done(pe_40_done)
  );
  
  std_reg #(32) down_34_write (
      .in(down_34_write_in),
      .write_en(down_34_write_write_en),
      .clk(clk),
      .out(down_34_write_out),
      .done(down_34_write_done)
  );
  
  std_reg #(32) left_34_read (
      .in(left_34_read_in),
      .write_en(left_34_read_write_en),
      .clk(clk),
      .out(left_34_read_out),
      .done(left_34_read_done)
  );
  
  std_reg #(32) top_34_read (
      .in(top_34_read_in),
      .write_en(top_34_read_write_en),
      .clk(clk),
      .out(top_34_read_out),
      .done(top_34_read_done)
  );
  
  mac_pe #() pe_34 (
      .top(pe_34_top),
      .left(pe_34_left),
      .go(pe_34_go),
      .clk(clk),
      .down(pe_34_down),
      .right(pe_34_right),
      .out(pe_34_out),
      .done(pe_34_done)
  );
  
  std_reg #(32) down_33_write (
      .in(down_33_write_in),
      .write_en(down_33_write_write_en),
      .clk(clk),
      .out(down_33_write_out),
      .done(down_33_write_done)
  );
  
  std_reg #(32) right_33_write (
      .in(right_33_write_in),
      .write_en(right_33_write_write_en),
      .clk(clk),
      .out(right_33_write_out),
      .done(right_33_write_done)
  );
  
  std_reg #(32) left_33_read (
      .in(left_33_read_in),
      .write_en(left_33_read_write_en),
      .clk(clk),
      .out(left_33_read_out),
      .done(left_33_read_done)
  );
  
  std_reg #(32) top_33_read (
      .in(top_33_read_in),
      .write_en(top_33_read_write_en),
      .clk(clk),
      .out(top_33_read_out),
      .done(top_33_read_done)
  );
  
  mac_pe #() pe_33 (
      .top(pe_33_top),
      .left(pe_33_left),
      .go(pe_33_go),
      .clk(clk),
      .down(pe_33_down),
      .right(pe_33_right),
      .out(pe_33_out),
      .done(pe_33_done)
  );
  
  std_reg #(32) down_32_write (
      .in(down_32_write_in),
      .write_en(down_32_write_write_en),
      .clk(clk),
      .out(down_32_write_out),
      .done(down_32_write_done)
  );
  
  std_reg #(32) right_32_write (
      .in(right_32_write_in),
      .write_en(right_32_write_write_en),
      .clk(clk),
      .out(right_32_write_out),
      .done(right_32_write_done)
  );
  
  std_reg #(32) left_32_read (
      .in(left_32_read_in),
      .write_en(left_32_read_write_en),
      .clk(clk),
      .out(left_32_read_out),
      .done(left_32_read_done)
  );
  
  std_reg #(32) top_32_read (
      .in(top_32_read_in),
      .write_en(top_32_read_write_en),
      .clk(clk),
      .out(top_32_read_out),
      .done(top_32_read_done)
  );
  
  mac_pe #() pe_32 (
      .top(pe_32_top),
      .left(pe_32_left),
      .go(pe_32_go),
      .clk(clk),
      .down(pe_32_down),
      .right(pe_32_right),
      .out(pe_32_out),
      .done(pe_32_done)
  );
  
  std_reg #(32) down_31_write (
      .in(down_31_write_in),
      .write_en(down_31_write_write_en),
      .clk(clk),
      .out(down_31_write_out),
      .done(down_31_write_done)
  );
  
  std_reg #(32) right_31_write (
      .in(right_31_write_in),
      .write_en(right_31_write_write_en),
      .clk(clk),
      .out(right_31_write_out),
      .done(right_31_write_done)
  );
  
  std_reg #(32) left_31_read (
      .in(left_31_read_in),
      .write_en(left_31_read_write_en),
      .clk(clk),
      .out(left_31_read_out),
      .done(left_31_read_done)
  );
  
  std_reg #(32) top_31_read (
      .in(top_31_read_in),
      .write_en(top_31_read_write_en),
      .clk(clk),
      .out(top_31_read_out),
      .done(top_31_read_done)
  );
  
  mac_pe #() pe_31 (
      .top(pe_31_top),
      .left(pe_31_left),
      .go(pe_31_go),
      .clk(clk),
      .down(pe_31_down),
      .right(pe_31_right),
      .out(pe_31_out),
      .done(pe_31_done)
  );
  
  std_reg #(32) down_30_write (
      .in(down_30_write_in),
      .write_en(down_30_write_write_en),
      .clk(clk),
      .out(down_30_write_out),
      .done(down_30_write_done)
  );
  
  std_reg #(32) right_30_write (
      .in(right_30_write_in),
      .write_en(right_30_write_write_en),
      .clk(clk),
      .out(right_30_write_out),
      .done(right_30_write_done)
  );
  
  std_reg #(32) left_30_read (
      .in(left_30_read_in),
      .write_en(left_30_read_write_en),
      .clk(clk),
      .out(left_30_read_out),
      .done(left_30_read_done)
  );
  
  std_reg #(32) top_30_read (
      .in(top_30_read_in),
      .write_en(top_30_read_write_en),
      .clk(clk),
      .out(top_30_read_out),
      .done(top_30_read_done)
  );
  
  mac_pe #() pe_30 (
      .top(pe_30_top),
      .left(pe_30_left),
      .go(pe_30_go),
      .clk(clk),
      .down(pe_30_down),
      .right(pe_30_right),
      .out(pe_30_out),
      .done(pe_30_done)
  );
  
  std_reg #(32) down_24_write (
      .in(down_24_write_in),
      .write_en(down_24_write_write_en),
      .clk(clk),
      .out(down_24_write_out),
      .done(down_24_write_done)
  );
  
  std_reg #(32) left_24_read (
      .in(left_24_read_in),
      .write_en(left_24_read_write_en),
      .clk(clk),
      .out(left_24_read_out),
      .done(left_24_read_done)
  );
  
  std_reg #(32) top_24_read (
      .in(top_24_read_in),
      .write_en(top_24_read_write_en),
      .clk(clk),
      .out(top_24_read_out),
      .done(top_24_read_done)
  );
  
  mac_pe #() pe_24 (
      .top(pe_24_top),
      .left(pe_24_left),
      .go(pe_24_go),
      .clk(clk),
      .down(pe_24_down),
      .right(pe_24_right),
      .out(pe_24_out),
      .done(pe_24_done)
  );
  
  std_reg #(32) down_23_write (
      .in(down_23_write_in),
      .write_en(down_23_write_write_en),
      .clk(clk),
      .out(down_23_write_out),
      .done(down_23_write_done)
  );
  
  std_reg #(32) right_23_write (
      .in(right_23_write_in),
      .write_en(right_23_write_write_en),
      .clk(clk),
      .out(right_23_write_out),
      .done(right_23_write_done)
  );
  
  std_reg #(32) left_23_read (
      .in(left_23_read_in),
      .write_en(left_23_read_write_en),
      .clk(clk),
      .out(left_23_read_out),
      .done(left_23_read_done)
  );
  
  std_reg #(32) top_23_read (
      .in(top_23_read_in),
      .write_en(top_23_read_write_en),
      .clk(clk),
      .out(top_23_read_out),
      .done(top_23_read_done)
  );
  
  mac_pe #() pe_23 (
      .top(pe_23_top),
      .left(pe_23_left),
      .go(pe_23_go),
      .clk(clk),
      .down(pe_23_down),
      .right(pe_23_right),
      .out(pe_23_out),
      .done(pe_23_done)
  );
  
  std_reg #(32) down_22_write (
      .in(down_22_write_in),
      .write_en(down_22_write_write_en),
      .clk(clk),
      .out(down_22_write_out),
      .done(down_22_write_done)
  );
  
  std_reg #(32) right_22_write (
      .in(right_22_write_in),
      .write_en(right_22_write_write_en),
      .clk(clk),
      .out(right_22_write_out),
      .done(right_22_write_done)
  );
  
  std_reg #(32) left_22_read (
      .in(left_22_read_in),
      .write_en(left_22_read_write_en),
      .clk(clk),
      .out(left_22_read_out),
      .done(left_22_read_done)
  );
  
  std_reg #(32) top_22_read (
      .in(top_22_read_in),
      .write_en(top_22_read_write_en),
      .clk(clk),
      .out(top_22_read_out),
      .done(top_22_read_done)
  );
  
  mac_pe #() pe_22 (
      .top(pe_22_top),
      .left(pe_22_left),
      .go(pe_22_go),
      .clk(clk),
      .down(pe_22_down),
      .right(pe_22_right),
      .out(pe_22_out),
      .done(pe_22_done)
  );
  
  std_reg #(32) down_21_write (
      .in(down_21_write_in),
      .write_en(down_21_write_write_en),
      .clk(clk),
      .out(down_21_write_out),
      .done(down_21_write_done)
  );
  
  std_reg #(32) right_21_write (
      .in(right_21_write_in),
      .write_en(right_21_write_write_en),
      .clk(clk),
      .out(right_21_write_out),
      .done(right_21_write_done)
  );
  
  std_reg #(32) left_21_read (
      .in(left_21_read_in),
      .write_en(left_21_read_write_en),
      .clk(clk),
      .out(left_21_read_out),
      .done(left_21_read_done)
  );
  
  std_reg #(32) top_21_read (
      .in(top_21_read_in),
      .write_en(top_21_read_write_en),
      .clk(clk),
      .out(top_21_read_out),
      .done(top_21_read_done)
  );
  
  mac_pe #() pe_21 (
      .top(pe_21_top),
      .left(pe_21_left),
      .go(pe_21_go),
      .clk(clk),
      .down(pe_21_down),
      .right(pe_21_right),
      .out(pe_21_out),
      .done(pe_21_done)
  );
  
  std_reg #(32) down_20_write (
      .in(down_20_write_in),
      .write_en(down_20_write_write_en),
      .clk(clk),
      .out(down_20_write_out),
      .done(down_20_write_done)
  );
  
  std_reg #(32) right_20_write (
      .in(right_20_write_in),
      .write_en(right_20_write_write_en),
      .clk(clk),
      .out(right_20_write_out),
      .done(right_20_write_done)
  );
  
  std_reg #(32) left_20_read (
      .in(left_20_read_in),
      .write_en(left_20_read_write_en),
      .clk(clk),
      .out(left_20_read_out),
      .done(left_20_read_done)
  );
  
  std_reg #(32) top_20_read (
      .in(top_20_read_in),
      .write_en(top_20_read_write_en),
      .clk(clk),
      .out(top_20_read_out),
      .done(top_20_read_done)
  );
  
  mac_pe #() pe_20 (
      .top(pe_20_top),
      .left(pe_20_left),
      .go(pe_20_go),
      .clk(clk),
      .down(pe_20_down),
      .right(pe_20_right),
      .out(pe_20_out),
      .done(pe_20_done)
  );
  
  std_reg #(32) down_14_write (
      .in(down_14_write_in),
      .write_en(down_14_write_write_en),
      .clk(clk),
      .out(down_14_write_out),
      .done(down_14_write_done)
  );
  
  std_reg #(32) left_14_read (
      .in(left_14_read_in),
      .write_en(left_14_read_write_en),
      .clk(clk),
      .out(left_14_read_out),
      .done(left_14_read_done)
  );
  
  std_reg #(32) top_14_read (
      .in(top_14_read_in),
      .write_en(top_14_read_write_en),
      .clk(clk),
      .out(top_14_read_out),
      .done(top_14_read_done)
  );
  
  mac_pe #() pe_14 (
      .top(pe_14_top),
      .left(pe_14_left),
      .go(pe_14_go),
      .clk(clk),
      .down(pe_14_down),
      .right(pe_14_right),
      .out(pe_14_out),
      .done(pe_14_done)
  );
  
  std_reg #(32) down_13_write (
      .in(down_13_write_in),
      .write_en(down_13_write_write_en),
      .clk(clk),
      .out(down_13_write_out),
      .done(down_13_write_done)
  );
  
  std_reg #(32) right_13_write (
      .in(right_13_write_in),
      .write_en(right_13_write_write_en),
      .clk(clk),
      .out(right_13_write_out),
      .done(right_13_write_done)
  );
  
  std_reg #(32) left_13_read (
      .in(left_13_read_in),
      .write_en(left_13_read_write_en),
      .clk(clk),
      .out(left_13_read_out),
      .done(left_13_read_done)
  );
  
  std_reg #(32) top_13_read (
      .in(top_13_read_in),
      .write_en(top_13_read_write_en),
      .clk(clk),
      .out(top_13_read_out),
      .done(top_13_read_done)
  );
  
  mac_pe #() pe_13 (
      .top(pe_13_top),
      .left(pe_13_left),
      .go(pe_13_go),
      .clk(clk),
      .down(pe_13_down),
      .right(pe_13_right),
      .out(pe_13_out),
      .done(pe_13_done)
  );
  
  std_reg #(32) down_12_write (
      .in(down_12_write_in),
      .write_en(down_12_write_write_en),
      .clk(clk),
      .out(down_12_write_out),
      .done(down_12_write_done)
  );
  
  std_reg #(32) right_12_write (
      .in(right_12_write_in),
      .write_en(right_12_write_write_en),
      .clk(clk),
      .out(right_12_write_out),
      .done(right_12_write_done)
  );
  
  std_reg #(32) left_12_read (
      .in(left_12_read_in),
      .write_en(left_12_read_write_en),
      .clk(clk),
      .out(left_12_read_out),
      .done(left_12_read_done)
  );
  
  std_reg #(32) top_12_read (
      .in(top_12_read_in),
      .write_en(top_12_read_write_en),
      .clk(clk),
      .out(top_12_read_out),
      .done(top_12_read_done)
  );
  
  mac_pe #() pe_12 (
      .top(pe_12_top),
      .left(pe_12_left),
      .go(pe_12_go),
      .clk(clk),
      .down(pe_12_down),
      .right(pe_12_right),
      .out(pe_12_out),
      .done(pe_12_done)
  );
  
  std_reg #(32) down_11_write (
      .in(down_11_write_in),
      .write_en(down_11_write_write_en),
      .clk(clk),
      .out(down_11_write_out),
      .done(down_11_write_done)
  );
  
  std_reg #(32) right_11_write (
      .in(right_11_write_in),
      .write_en(right_11_write_write_en),
      .clk(clk),
      .out(right_11_write_out),
      .done(right_11_write_done)
  );
  
  std_reg #(32) left_11_read (
      .in(left_11_read_in),
      .write_en(left_11_read_write_en),
      .clk(clk),
      .out(left_11_read_out),
      .done(left_11_read_done)
  );
  
  std_reg #(32) top_11_read (
      .in(top_11_read_in),
      .write_en(top_11_read_write_en),
      .clk(clk),
      .out(top_11_read_out),
      .done(top_11_read_done)
  );
  
  mac_pe #() pe_11 (
      .top(pe_11_top),
      .left(pe_11_left),
      .go(pe_11_go),
      .clk(clk),
      .down(pe_11_down),
      .right(pe_11_right),
      .out(pe_11_out),
      .done(pe_11_done)
  );
  
  std_reg #(32) down_10_write (
      .in(down_10_write_in),
      .write_en(down_10_write_write_en),
      .clk(clk),
      .out(down_10_write_out),
      .done(down_10_write_done)
  );
  
  std_reg #(32) right_10_write (
      .in(right_10_write_in),
      .write_en(right_10_write_write_en),
      .clk(clk),
      .out(right_10_write_out),
      .done(right_10_write_done)
  );
  
  std_reg #(32) left_10_read (
      .in(left_10_read_in),
      .write_en(left_10_read_write_en),
      .clk(clk),
      .out(left_10_read_out),
      .done(left_10_read_done)
  );
  
  std_reg #(32) top_10_read (
      .in(top_10_read_in),
      .write_en(top_10_read_write_en),
      .clk(clk),
      .out(top_10_read_out),
      .done(top_10_read_done)
  );
  
  mac_pe #() pe_10 (
      .top(pe_10_top),
      .left(pe_10_left),
      .go(pe_10_go),
      .clk(clk),
      .down(pe_10_down),
      .right(pe_10_right),
      .out(pe_10_out),
      .done(pe_10_done)
  );
  
  std_reg #(32) down_04_write (
      .in(down_04_write_in),
      .write_en(down_04_write_write_en),
      .clk(clk),
      .out(down_04_write_out),
      .done(down_04_write_done)
  );
  
  std_reg #(32) left_04_read (
      .in(left_04_read_in),
      .write_en(left_04_read_write_en),
      .clk(clk),
      .out(left_04_read_out),
      .done(left_04_read_done)
  );
  
  std_reg #(32) top_04_read (
      .in(top_04_read_in),
      .write_en(top_04_read_write_en),
      .clk(clk),
      .out(top_04_read_out),
      .done(top_04_read_done)
  );
  
  mac_pe #() pe_04 (
      .top(pe_04_top),
      .left(pe_04_left),
      .go(pe_04_go),
      .clk(clk),
      .down(pe_04_down),
      .right(pe_04_right),
      .out(pe_04_out),
      .done(pe_04_done)
  );
  
  std_reg #(32) down_03_write (
      .in(down_03_write_in),
      .write_en(down_03_write_write_en),
      .clk(clk),
      .out(down_03_write_out),
      .done(down_03_write_done)
  );
  
  std_reg #(32) right_03_write (
      .in(right_03_write_in),
      .write_en(right_03_write_write_en),
      .clk(clk),
      .out(right_03_write_out),
      .done(right_03_write_done)
  );
  
  std_reg #(32) left_03_read (
      .in(left_03_read_in),
      .write_en(left_03_read_write_en),
      .clk(clk),
      .out(left_03_read_out),
      .done(left_03_read_done)
  );
  
  std_reg #(32) top_03_read (
      .in(top_03_read_in),
      .write_en(top_03_read_write_en),
      .clk(clk),
      .out(top_03_read_out),
      .done(top_03_read_done)
  );
  
  mac_pe #() pe_03 (
      .top(pe_03_top),
      .left(pe_03_left),
      .go(pe_03_go),
      .clk(clk),
      .down(pe_03_down),
      .right(pe_03_right),
      .out(pe_03_out),
      .done(pe_03_done)
  );
  
  std_reg #(32) down_02_write (
      .in(down_02_write_in),
      .write_en(down_02_write_write_en),
      .clk(clk),
      .out(down_02_write_out),
      .done(down_02_write_done)
  );
  
  std_reg #(32) right_02_write (
      .in(right_02_write_in),
      .write_en(right_02_write_write_en),
      .clk(clk),
      .out(right_02_write_out),
      .done(right_02_write_done)
  );
  
  std_reg #(32) left_02_read (
      .in(left_02_read_in),
      .write_en(left_02_read_write_en),
      .clk(clk),
      .out(left_02_read_out),
      .done(left_02_read_done)
  );
  
  std_reg #(32) top_02_read (
      .in(top_02_read_in),
      .write_en(top_02_read_write_en),
      .clk(clk),
      .out(top_02_read_out),
      .done(top_02_read_done)
  );
  
  mac_pe #() pe_02 (
      .top(pe_02_top),
      .left(pe_02_left),
      .go(pe_02_go),
      .clk(clk),
      .down(pe_02_down),
      .right(pe_02_right),
      .out(pe_02_out),
      .done(pe_02_done)
  );
  
  std_reg #(32) down_01_write (
      .in(down_01_write_in),
      .write_en(down_01_write_write_en),
      .clk(clk),
      .out(down_01_write_out),
      .done(down_01_write_done)
  );
  
  std_reg #(32) right_01_write (
      .in(right_01_write_in),
      .write_en(right_01_write_write_en),
      .clk(clk),
      .out(right_01_write_out),
      .done(right_01_write_done)
  );
  
  std_reg #(32) left_01_read (
      .in(left_01_read_in),
      .write_en(left_01_read_write_en),
      .clk(clk),
      .out(left_01_read_out),
      .done(left_01_read_done)
  );
  
  std_reg #(32) top_01_read (
      .in(top_01_read_in),
      .write_en(top_01_read_write_en),
      .clk(clk),
      .out(top_01_read_out),
      .done(top_01_read_done)
  );
  
  mac_pe #() pe_01 (
      .top(pe_01_top),
      .left(pe_01_left),
      .go(pe_01_go),
      .clk(clk),
      .down(pe_01_down),
      .right(pe_01_right),
      .out(pe_01_out),
      .done(pe_01_done)
  );
  
  std_reg #(32) down_00_write (
      .in(down_00_write_in),
      .write_en(down_00_write_write_en),
      .clk(clk),
      .out(down_00_write_out),
      .done(down_00_write_done)
  );
  
  std_reg #(32) right_00_write (
      .in(right_00_write_in),
      .write_en(right_00_write_write_en),
      .clk(clk),
      .out(right_00_write_out),
      .done(right_00_write_done)
  );
  
  std_reg #(32) left_00_read (
      .in(left_00_read_in),
      .write_en(left_00_read_write_en),
      .clk(clk),
      .out(left_00_read_out),
      .done(left_00_read_done)
  );
  
  std_reg #(32) top_00_read (
      .in(top_00_read_in),
      .write_en(top_00_read_write_en),
      .clk(clk),
      .out(top_00_read_out),
      .done(top_00_read_done)
  );
  
  mac_pe #() pe_00 (
      .top(pe_00_top),
      .left(pe_00_left),
      .go(pe_00_go),
      .clk(clk),
      .down(pe_00_down),
      .right(pe_00_right),
      .out(pe_00_out),
      .done(pe_00_done)
  );
  
  std_mem_d1 #(32, 5, 3) l4 (
      .addr0(l4_addr0),
      .write_data(l4_write_data),
      .write_en(l4_write_en),
      .clk(clk),
      .read_data(l4_read_data),
      .done(l4_done)
  );
  
  std_add #(3) l4_add (
      .left(l4_add_left),
      .right(l4_add_right),
      .out(l4_add_out)
  );
  
  std_reg #(3) l4_idx (
      .in(l4_idx_in),
      .write_en(l4_idx_write_en),
      .clk(clk),
      .out(l4_idx_out),
      .done(l4_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) l3 (
      .addr0(l3_addr0),
      .write_data(l3_write_data),
      .write_en(l3_write_en),
      .clk(clk),
      .read_data(l3_read_data),
      .done(l3_done)
  );
  
  std_add #(3) l3_add (
      .left(l3_add_left),
      .right(l3_add_right),
      .out(l3_add_out)
  );
  
  std_reg #(3) l3_idx (
      .in(l3_idx_in),
      .write_en(l3_idx_write_en),
      .clk(clk),
      .out(l3_idx_out),
      .done(l3_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) l2 (
      .addr0(l2_addr0),
      .write_data(l2_write_data),
      .write_en(l2_write_en),
      .clk(clk),
      .read_data(l2_read_data),
      .done(l2_done)
  );
  
  std_add #(3) l2_add (
      .left(l2_add_left),
      .right(l2_add_right),
      .out(l2_add_out)
  );
  
  std_reg #(3) l2_idx (
      .in(l2_idx_in),
      .write_en(l2_idx_write_en),
      .clk(clk),
      .out(l2_idx_out),
      .done(l2_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) l1 (
      .addr0(l1_addr0),
      .write_data(l1_write_data),
      .write_en(l1_write_en),
      .clk(clk),
      .read_data(l1_read_data),
      .done(l1_done)
  );
  
  std_add #(3) l1_add (
      .left(l1_add_left),
      .right(l1_add_right),
      .out(l1_add_out)
  );
  
  std_reg #(3) l1_idx (
      .in(l1_idx_in),
      .write_en(l1_idx_write_en),
      .clk(clk),
      .out(l1_idx_out),
      .done(l1_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) l0 (
      .addr0(l0_addr0),
      .write_data(l0_write_data),
      .write_en(l0_write_en),
      .clk(clk),
      .read_data(l0_read_data),
      .done(l0_done)
  );
  
  std_add #(3) l0_add (
      .left(l0_add_left),
      .right(l0_add_right),
      .out(l0_add_out)
  );
  
  std_reg #(3) l0_idx (
      .in(l0_idx_in),
      .write_en(l0_idx_write_en),
      .clk(clk),
      .out(l0_idx_out),
      .done(l0_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) t4 (
      .addr0(t4_addr0),
      .write_data(t4_write_data),
      .write_en(t4_write_en),
      .clk(clk),
      .read_data(t4_read_data),
      .done(t4_done)
  );
  
  std_add #(3) t4_add (
      .left(t4_add_left),
      .right(t4_add_right),
      .out(t4_add_out)
  );
  
  std_reg #(3) t4_idx (
      .in(t4_idx_in),
      .write_en(t4_idx_write_en),
      .clk(clk),
      .out(t4_idx_out),
      .done(t4_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) t3 (
      .addr0(t3_addr0),
      .write_data(t3_write_data),
      .write_en(t3_write_en),
      .clk(clk),
      .read_data(t3_read_data),
      .done(t3_done)
  );
  
  std_add #(3) t3_add (
      .left(t3_add_left),
      .right(t3_add_right),
      .out(t3_add_out)
  );
  
  std_reg #(3) t3_idx (
      .in(t3_idx_in),
      .write_en(t3_idx_write_en),
      .clk(clk),
      .out(t3_idx_out),
      .done(t3_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) t2 (
      .addr0(t2_addr0),
      .write_data(t2_write_data),
      .write_en(t2_write_en),
      .clk(clk),
      .read_data(t2_read_data),
      .done(t2_done)
  );
  
  std_add #(3) t2_add (
      .left(t2_add_left),
      .right(t2_add_right),
      .out(t2_add_out)
  );
  
  std_reg #(3) t2_idx (
      .in(t2_idx_in),
      .write_en(t2_idx_write_en),
      .clk(clk),
      .out(t2_idx_out),
      .done(t2_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) t1 (
      .addr0(t1_addr0),
      .write_data(t1_write_data),
      .write_en(t1_write_en),
      .clk(clk),
      .read_data(t1_read_data),
      .done(t1_done)
  );
  
  std_add #(3) t1_add (
      .left(t1_add_left),
      .right(t1_add_right),
      .out(t1_add_out)
  );
  
  std_reg #(3) t1_idx (
      .in(t1_idx_in),
      .write_en(t1_idx_write_en),
      .clk(clk),
      .out(t1_idx_out),
      .done(t1_idx_done)
  );
  
  std_mem_d1 #(32, 5, 3) t0 (
      .addr0(t0_addr0),
      .write_data(t0_write_data),
      .write_en(t0_write_en),
      .clk(clk),
      .read_data(t0_read_data),
      .done(t0_done)
  );
  
  std_add #(3) t0_add (
      .left(t0_add_left),
      .right(t0_add_right),
      .out(t0_add_out)
  );
  
  std_reg #(3) t0_idx (
      .in(t0_idx_in),
      .write_en(t0_idx_write_en),
      .clk(clk),
      .out(t0_idx_out),
      .done(t0_idx_done)
  );
  
  std_reg #(1) par_reset0 (
      .in(par_reset0_in),
      .write_en(par_reset0_write_en),
      .clk(clk),
      .out(par_reset0_out),
      .done(par_reset0_done)
  );
  
  std_reg #(1) par_done_reg0 (
      .in(par_done_reg0_in),
      .write_en(par_done_reg0_write_en),
      .clk(clk),
      .out(par_done_reg0_out),
      .done(par_done_reg0_done)
  );
  
  std_reg #(1) par_done_reg1 (
      .in(par_done_reg1_in),
      .write_en(par_done_reg1_write_en),
      .clk(clk),
      .out(par_done_reg1_out),
      .done(par_done_reg1_done)
  );
  
  std_reg #(1) par_done_reg2 (
      .in(par_done_reg2_in),
      .write_en(par_done_reg2_write_en),
      .clk(clk),
      .out(par_done_reg2_out),
      .done(par_done_reg2_done)
  );
  
  std_reg #(1) par_done_reg3 (
      .in(par_done_reg3_in),
      .write_en(par_done_reg3_write_en),
      .clk(clk),
      .out(par_done_reg3_out),
      .done(par_done_reg3_done)
  );
  
  std_reg #(1) par_done_reg4 (
      .in(par_done_reg4_in),
      .write_en(par_done_reg4_write_en),
      .clk(clk),
      .out(par_done_reg4_out),
      .done(par_done_reg4_done)
  );
  
  std_reg #(1) par_done_reg5 (
      .in(par_done_reg5_in),
      .write_en(par_done_reg5_write_en),
      .clk(clk),
      .out(par_done_reg5_out),
      .done(par_done_reg5_done)
  );
  
  std_reg #(1) par_done_reg6 (
      .in(par_done_reg6_in),
      .write_en(par_done_reg6_write_en),
      .clk(clk),
      .out(par_done_reg6_out),
      .done(par_done_reg6_done)
  );
  
  std_reg #(1) par_done_reg7 (
      .in(par_done_reg7_in),
      .write_en(par_done_reg7_write_en),
      .clk(clk),
      .out(par_done_reg7_out),
      .done(par_done_reg7_done)
  );
  
  std_reg #(1) par_done_reg8 (
      .in(par_done_reg8_in),
      .write_en(par_done_reg8_write_en),
      .clk(clk),
      .out(par_done_reg8_out),
      .done(par_done_reg8_done)
  );
  
  std_reg #(1) par_done_reg9 (
      .in(par_done_reg9_in),
      .write_en(par_done_reg9_write_en),
      .clk(clk),
      .out(par_done_reg9_out),
      .done(par_done_reg9_done)
  );
  
  std_reg #(1) par_reset1 (
      .in(par_reset1_in),
      .write_en(par_reset1_write_en),
      .clk(clk),
      .out(par_reset1_out),
      .done(par_reset1_done)
  );
  
  std_reg #(1) par_done_reg10 (
      .in(par_done_reg10_in),
      .write_en(par_done_reg10_write_en),
      .clk(clk),
      .out(par_done_reg10_out),
      .done(par_done_reg10_done)
  );
  
  std_reg #(1) par_done_reg11 (
      .in(par_done_reg11_in),
      .write_en(par_done_reg11_write_en),
      .clk(clk),
      .out(par_done_reg11_out),
      .done(par_done_reg11_done)
  );
  
  std_reg #(1) par_reset2 (
      .in(par_reset2_in),
      .write_en(par_reset2_write_en),
      .clk(clk),
      .out(par_reset2_out),
      .done(par_reset2_done)
  );
  
  std_reg #(1) par_done_reg12 (
      .in(par_done_reg12_in),
      .write_en(par_done_reg12_write_en),
      .clk(clk),
      .out(par_done_reg12_out),
      .done(par_done_reg12_done)
  );
  
  std_reg #(1) par_done_reg13 (
      .in(par_done_reg13_in),
      .write_en(par_done_reg13_write_en),
      .clk(clk),
      .out(par_done_reg13_out),
      .done(par_done_reg13_done)
  );
  
  std_reg #(1) par_reset3 (
      .in(par_reset3_in),
      .write_en(par_reset3_write_en),
      .clk(clk),
      .out(par_reset3_out),
      .done(par_reset3_done)
  );
  
  std_reg #(1) par_done_reg14 (
      .in(par_done_reg14_in),
      .write_en(par_done_reg14_write_en),
      .clk(clk),
      .out(par_done_reg14_out),
      .done(par_done_reg14_done)
  );
  
  std_reg #(1) par_done_reg15 (
      .in(par_done_reg15_in),
      .write_en(par_done_reg15_write_en),
      .clk(clk),
      .out(par_done_reg15_out),
      .done(par_done_reg15_done)
  );
  
  std_reg #(1) par_done_reg16 (
      .in(par_done_reg16_in),
      .write_en(par_done_reg16_write_en),
      .clk(clk),
      .out(par_done_reg16_out),
      .done(par_done_reg16_done)
  );
  
  std_reg #(1) par_done_reg17 (
      .in(par_done_reg17_in),
      .write_en(par_done_reg17_write_en),
      .clk(clk),
      .out(par_done_reg17_out),
      .done(par_done_reg17_done)
  );
  
  std_reg #(1) par_done_reg18 (
      .in(par_done_reg18_in),
      .write_en(par_done_reg18_write_en),
      .clk(clk),
      .out(par_done_reg18_out),
      .done(par_done_reg18_done)
  );
  
  std_reg #(1) par_reset4 (
      .in(par_reset4_in),
      .write_en(par_reset4_write_en),
      .clk(clk),
      .out(par_reset4_out),
      .done(par_reset4_done)
  );
  
  std_reg #(1) par_done_reg19 (
      .in(par_done_reg19_in),
      .write_en(par_done_reg19_write_en),
      .clk(clk),
      .out(par_done_reg19_out),
      .done(par_done_reg19_done)
  );
  
  std_reg #(1) par_done_reg20 (
      .in(par_done_reg20_in),
      .write_en(par_done_reg20_write_en),
      .clk(clk),
      .out(par_done_reg20_out),
      .done(par_done_reg20_done)
  );
  
  std_reg #(1) par_done_reg21 (
      .in(par_done_reg21_in),
      .write_en(par_done_reg21_write_en),
      .clk(clk),
      .out(par_done_reg21_out),
      .done(par_done_reg21_done)
  );
  
  std_reg #(1) par_done_reg22 (
      .in(par_done_reg22_in),
      .write_en(par_done_reg22_write_en),
      .clk(clk),
      .out(par_done_reg22_out),
      .done(par_done_reg22_done)
  );
  
  std_reg #(1) par_done_reg23 (
      .in(par_done_reg23_in),
      .write_en(par_done_reg23_write_en),
      .clk(clk),
      .out(par_done_reg23_out),
      .done(par_done_reg23_done)
  );
  
  std_reg #(1) par_done_reg24 (
      .in(par_done_reg24_in),
      .write_en(par_done_reg24_write_en),
      .clk(clk),
      .out(par_done_reg24_out),
      .done(par_done_reg24_done)
  );
  
  std_reg #(1) par_reset5 (
      .in(par_reset5_in),
      .write_en(par_reset5_write_en),
      .clk(clk),
      .out(par_reset5_out),
      .done(par_reset5_done)
  );
  
  std_reg #(1) par_done_reg25 (
      .in(par_done_reg25_in),
      .write_en(par_done_reg25_write_en),
      .clk(clk),
      .out(par_done_reg25_out),
      .done(par_done_reg25_done)
  );
  
  std_reg #(1) par_done_reg26 (
      .in(par_done_reg26_in),
      .write_en(par_done_reg26_write_en),
      .clk(clk),
      .out(par_done_reg26_out),
      .done(par_done_reg26_done)
  );
  
  std_reg #(1) par_done_reg27 (
      .in(par_done_reg27_in),
      .write_en(par_done_reg27_write_en),
      .clk(clk),
      .out(par_done_reg27_out),
      .done(par_done_reg27_done)
  );
  
  std_reg #(1) par_done_reg28 (
      .in(par_done_reg28_in),
      .write_en(par_done_reg28_write_en),
      .clk(clk),
      .out(par_done_reg28_out),
      .done(par_done_reg28_done)
  );
  
  std_reg #(1) par_done_reg29 (
      .in(par_done_reg29_in),
      .write_en(par_done_reg29_write_en),
      .clk(clk),
      .out(par_done_reg29_out),
      .done(par_done_reg29_done)
  );
  
  std_reg #(1) par_done_reg30 (
      .in(par_done_reg30_in),
      .write_en(par_done_reg30_write_en),
      .clk(clk),
      .out(par_done_reg30_out),
      .done(par_done_reg30_done)
  );
  
  std_reg #(1) par_done_reg31 (
      .in(par_done_reg31_in),
      .write_en(par_done_reg31_write_en),
      .clk(clk),
      .out(par_done_reg31_out),
      .done(par_done_reg31_done)
  );
  
  std_reg #(1) par_done_reg32 (
      .in(par_done_reg32_in),
      .write_en(par_done_reg32_write_en),
      .clk(clk),
      .out(par_done_reg32_out),
      .done(par_done_reg32_done)
  );
  
  std_reg #(1) par_done_reg33 (
      .in(par_done_reg33_in),
      .write_en(par_done_reg33_write_en),
      .clk(clk),
      .out(par_done_reg33_out),
      .done(par_done_reg33_done)
  );
  
  std_reg #(1) par_reset6 (
      .in(par_reset6_in),
      .write_en(par_reset6_write_en),
      .clk(clk),
      .out(par_reset6_out),
      .done(par_reset6_done)
  );
  
  std_reg #(1) par_done_reg34 (
      .in(par_done_reg34_in),
      .write_en(par_done_reg34_write_en),
      .clk(clk),
      .out(par_done_reg34_out),
      .done(par_done_reg34_done)
  );
  
  std_reg #(1) par_done_reg35 (
      .in(par_done_reg35_in),
      .write_en(par_done_reg35_write_en),
      .clk(clk),
      .out(par_done_reg35_out),
      .done(par_done_reg35_done)
  );
  
  std_reg #(1) par_done_reg36 (
      .in(par_done_reg36_in),
      .write_en(par_done_reg36_write_en),
      .clk(clk),
      .out(par_done_reg36_out),
      .done(par_done_reg36_done)
  );
  
  std_reg #(1) par_done_reg37 (
      .in(par_done_reg37_in),
      .write_en(par_done_reg37_write_en),
      .clk(clk),
      .out(par_done_reg37_out),
      .done(par_done_reg37_done)
  );
  
  std_reg #(1) par_done_reg38 (
      .in(par_done_reg38_in),
      .write_en(par_done_reg38_write_en),
      .clk(clk),
      .out(par_done_reg38_out),
      .done(par_done_reg38_done)
  );
  
  std_reg #(1) par_done_reg39 (
      .in(par_done_reg39_in),
      .write_en(par_done_reg39_write_en),
      .clk(clk),
      .out(par_done_reg39_out),
      .done(par_done_reg39_done)
  );
  
  std_reg #(1) par_done_reg40 (
      .in(par_done_reg40_in),
      .write_en(par_done_reg40_write_en),
      .clk(clk),
      .out(par_done_reg40_out),
      .done(par_done_reg40_done)
  );
  
  std_reg #(1) par_done_reg41 (
      .in(par_done_reg41_in),
      .write_en(par_done_reg41_write_en),
      .clk(clk),
      .out(par_done_reg41_out),
      .done(par_done_reg41_done)
  );
  
  std_reg #(1) par_done_reg42 (
      .in(par_done_reg42_in),
      .write_en(par_done_reg42_write_en),
      .clk(clk),
      .out(par_done_reg42_out),
      .done(par_done_reg42_done)
  );
  
  std_reg #(1) par_done_reg43 (
      .in(par_done_reg43_in),
      .write_en(par_done_reg43_write_en),
      .clk(clk),
      .out(par_done_reg43_out),
      .done(par_done_reg43_done)
  );
  
  std_reg #(1) par_done_reg44 (
      .in(par_done_reg44_in),
      .write_en(par_done_reg44_write_en),
      .clk(clk),
      .out(par_done_reg44_out),
      .done(par_done_reg44_done)
  );
  
  std_reg #(1) par_done_reg45 (
      .in(par_done_reg45_in),
      .write_en(par_done_reg45_write_en),
      .clk(clk),
      .out(par_done_reg45_out),
      .done(par_done_reg45_done)
  );
  
  std_reg #(1) par_reset7 (
      .in(par_reset7_in),
      .write_en(par_reset7_write_en),
      .clk(clk),
      .out(par_reset7_out),
      .done(par_reset7_done)
  );
  
  std_reg #(1) par_done_reg46 (
      .in(par_done_reg46_in),
      .write_en(par_done_reg46_write_en),
      .clk(clk),
      .out(par_done_reg46_out),
      .done(par_done_reg46_done)
  );
  
  std_reg #(1) par_done_reg47 (
      .in(par_done_reg47_in),
      .write_en(par_done_reg47_write_en),
      .clk(clk),
      .out(par_done_reg47_out),
      .done(par_done_reg47_done)
  );
  
  std_reg #(1) par_done_reg48 (
      .in(par_done_reg48_in),
      .write_en(par_done_reg48_write_en),
      .clk(clk),
      .out(par_done_reg48_out),
      .done(par_done_reg48_done)
  );
  
  std_reg #(1) par_done_reg49 (
      .in(par_done_reg49_in),
      .write_en(par_done_reg49_write_en),
      .clk(clk),
      .out(par_done_reg49_out),
      .done(par_done_reg49_done)
  );
  
  std_reg #(1) par_done_reg50 (
      .in(par_done_reg50_in),
      .write_en(par_done_reg50_write_en),
      .clk(clk),
      .out(par_done_reg50_out),
      .done(par_done_reg50_done)
  );
  
  std_reg #(1) par_done_reg51 (
      .in(par_done_reg51_in),
      .write_en(par_done_reg51_write_en),
      .clk(clk),
      .out(par_done_reg51_out),
      .done(par_done_reg51_done)
  );
  
  std_reg #(1) par_done_reg52 (
      .in(par_done_reg52_in),
      .write_en(par_done_reg52_write_en),
      .clk(clk),
      .out(par_done_reg52_out),
      .done(par_done_reg52_done)
  );
  
  std_reg #(1) par_done_reg53 (
      .in(par_done_reg53_in),
      .write_en(par_done_reg53_write_en),
      .clk(clk),
      .out(par_done_reg53_out),
      .done(par_done_reg53_done)
  );
  
  std_reg #(1) par_done_reg54 (
      .in(par_done_reg54_in),
      .write_en(par_done_reg54_write_en),
      .clk(clk),
      .out(par_done_reg54_out),
      .done(par_done_reg54_done)
  );
  
  std_reg #(1) par_done_reg55 (
      .in(par_done_reg55_in),
      .write_en(par_done_reg55_write_en),
      .clk(clk),
      .out(par_done_reg55_out),
      .done(par_done_reg55_done)
  );
  
  std_reg #(1) par_done_reg56 (
      .in(par_done_reg56_in),
      .write_en(par_done_reg56_write_en),
      .clk(clk),
      .out(par_done_reg56_out),
      .done(par_done_reg56_done)
  );
  
  std_reg #(1) par_done_reg57 (
      .in(par_done_reg57_in),
      .write_en(par_done_reg57_write_en),
      .clk(clk),
      .out(par_done_reg57_out),
      .done(par_done_reg57_done)
  );
  
  std_reg #(1) par_done_reg58 (
      .in(par_done_reg58_in),
      .write_en(par_done_reg58_write_en),
      .clk(clk),
      .out(par_done_reg58_out),
      .done(par_done_reg58_done)
  );
  
  std_reg #(1) par_done_reg59 (
      .in(par_done_reg59_in),
      .write_en(par_done_reg59_write_en),
      .clk(clk),
      .out(par_done_reg59_out),
      .done(par_done_reg59_done)
  );
  
  std_reg #(1) par_reset8 (
      .in(par_reset8_in),
      .write_en(par_reset8_write_en),
      .clk(clk),
      .out(par_reset8_out),
      .done(par_reset8_done)
  );
  
  std_reg #(1) par_done_reg60 (
      .in(par_done_reg60_in),
      .write_en(par_done_reg60_write_en),
      .clk(clk),
      .out(par_done_reg60_out),
      .done(par_done_reg60_done)
  );
  
  std_reg #(1) par_done_reg61 (
      .in(par_done_reg61_in),
      .write_en(par_done_reg61_write_en),
      .clk(clk),
      .out(par_done_reg61_out),
      .done(par_done_reg61_done)
  );
  
  std_reg #(1) par_done_reg62 (
      .in(par_done_reg62_in),
      .write_en(par_done_reg62_write_en),
      .clk(clk),
      .out(par_done_reg62_out),
      .done(par_done_reg62_done)
  );
  
  std_reg #(1) par_done_reg63 (
      .in(par_done_reg63_in),
      .write_en(par_done_reg63_write_en),
      .clk(clk),
      .out(par_done_reg63_out),
      .done(par_done_reg63_done)
  );
  
  std_reg #(1) par_done_reg64 (
      .in(par_done_reg64_in),
      .write_en(par_done_reg64_write_en),
      .clk(clk),
      .out(par_done_reg64_out),
      .done(par_done_reg64_done)
  );
  
  std_reg #(1) par_done_reg65 (
      .in(par_done_reg65_in),
      .write_en(par_done_reg65_write_en),
      .clk(clk),
      .out(par_done_reg65_out),
      .done(par_done_reg65_done)
  );
  
  std_reg #(1) par_done_reg66 (
      .in(par_done_reg66_in),
      .write_en(par_done_reg66_write_en),
      .clk(clk),
      .out(par_done_reg66_out),
      .done(par_done_reg66_done)
  );
  
  std_reg #(1) par_done_reg67 (
      .in(par_done_reg67_in),
      .write_en(par_done_reg67_write_en),
      .clk(clk),
      .out(par_done_reg67_out),
      .done(par_done_reg67_done)
  );
  
  std_reg #(1) par_done_reg68 (
      .in(par_done_reg68_in),
      .write_en(par_done_reg68_write_en),
      .clk(clk),
      .out(par_done_reg68_out),
      .done(par_done_reg68_done)
  );
  
  std_reg #(1) par_done_reg69 (
      .in(par_done_reg69_in),
      .write_en(par_done_reg69_write_en),
      .clk(clk),
      .out(par_done_reg69_out),
      .done(par_done_reg69_done)
  );
  
  std_reg #(1) par_done_reg70 (
      .in(par_done_reg70_in),
      .write_en(par_done_reg70_write_en),
      .clk(clk),
      .out(par_done_reg70_out),
      .done(par_done_reg70_done)
  );
  
  std_reg #(1) par_done_reg71 (
      .in(par_done_reg71_in),
      .write_en(par_done_reg71_write_en),
      .clk(clk),
      .out(par_done_reg71_out),
      .done(par_done_reg71_done)
  );
  
  std_reg #(1) par_done_reg72 (
      .in(par_done_reg72_in),
      .write_en(par_done_reg72_write_en),
      .clk(clk),
      .out(par_done_reg72_out),
      .done(par_done_reg72_done)
  );
  
  std_reg #(1) par_done_reg73 (
      .in(par_done_reg73_in),
      .write_en(par_done_reg73_write_en),
      .clk(clk),
      .out(par_done_reg73_out),
      .done(par_done_reg73_done)
  );
  
  std_reg #(1) par_done_reg74 (
      .in(par_done_reg74_in),
      .write_en(par_done_reg74_write_en),
      .clk(clk),
      .out(par_done_reg74_out),
      .done(par_done_reg74_done)
  );
  
  std_reg #(1) par_done_reg75 (
      .in(par_done_reg75_in),
      .write_en(par_done_reg75_write_en),
      .clk(clk),
      .out(par_done_reg75_out),
      .done(par_done_reg75_done)
  );
  
  std_reg #(1) par_done_reg76 (
      .in(par_done_reg76_in),
      .write_en(par_done_reg76_write_en),
      .clk(clk),
      .out(par_done_reg76_out),
      .done(par_done_reg76_done)
  );
  
  std_reg #(1) par_done_reg77 (
      .in(par_done_reg77_in),
      .write_en(par_done_reg77_write_en),
      .clk(clk),
      .out(par_done_reg77_out),
      .done(par_done_reg77_done)
  );
  
  std_reg #(1) par_done_reg78 (
      .in(par_done_reg78_in),
      .write_en(par_done_reg78_write_en),
      .clk(clk),
      .out(par_done_reg78_out),
      .done(par_done_reg78_done)
  );
  
  std_reg #(1) par_done_reg79 (
      .in(par_done_reg79_in),
      .write_en(par_done_reg79_write_en),
      .clk(clk),
      .out(par_done_reg79_out),
      .done(par_done_reg79_done)
  );
  
  std_reg #(1) par_reset9 (
      .in(par_reset9_in),
      .write_en(par_reset9_write_en),
      .clk(clk),
      .out(par_reset9_out),
      .done(par_reset9_done)
  );
  
  std_reg #(1) par_done_reg80 (
      .in(par_done_reg80_in),
      .write_en(par_done_reg80_write_en),
      .clk(clk),
      .out(par_done_reg80_out),
      .done(par_done_reg80_done)
  );
  
  std_reg #(1) par_done_reg81 (
      .in(par_done_reg81_in),
      .write_en(par_done_reg81_write_en),
      .clk(clk),
      .out(par_done_reg81_out),
      .done(par_done_reg81_done)
  );
  
  std_reg #(1) par_done_reg82 (
      .in(par_done_reg82_in),
      .write_en(par_done_reg82_write_en),
      .clk(clk),
      .out(par_done_reg82_out),
      .done(par_done_reg82_done)
  );
  
  std_reg #(1) par_done_reg83 (
      .in(par_done_reg83_in),
      .write_en(par_done_reg83_write_en),
      .clk(clk),
      .out(par_done_reg83_out),
      .done(par_done_reg83_done)
  );
  
  std_reg #(1) par_done_reg84 (
      .in(par_done_reg84_in),
      .write_en(par_done_reg84_write_en),
      .clk(clk),
      .out(par_done_reg84_out),
      .done(par_done_reg84_done)
  );
  
  std_reg #(1) par_done_reg85 (
      .in(par_done_reg85_in),
      .write_en(par_done_reg85_write_en),
      .clk(clk),
      .out(par_done_reg85_out),
      .done(par_done_reg85_done)
  );
  
  std_reg #(1) par_done_reg86 (
      .in(par_done_reg86_in),
      .write_en(par_done_reg86_write_en),
      .clk(clk),
      .out(par_done_reg86_out),
      .done(par_done_reg86_done)
  );
  
  std_reg #(1) par_done_reg87 (
      .in(par_done_reg87_in),
      .write_en(par_done_reg87_write_en),
      .clk(clk),
      .out(par_done_reg87_out),
      .done(par_done_reg87_done)
  );
  
  std_reg #(1) par_done_reg88 (
      .in(par_done_reg88_in),
      .write_en(par_done_reg88_write_en),
      .clk(clk),
      .out(par_done_reg88_out),
      .done(par_done_reg88_done)
  );
  
  std_reg #(1) par_done_reg89 (
      .in(par_done_reg89_in),
      .write_en(par_done_reg89_write_en),
      .clk(clk),
      .out(par_done_reg89_out),
      .done(par_done_reg89_done)
  );
  
  std_reg #(1) par_done_reg90 (
      .in(par_done_reg90_in),
      .write_en(par_done_reg90_write_en),
      .clk(clk),
      .out(par_done_reg90_out),
      .done(par_done_reg90_done)
  );
  
  std_reg #(1) par_done_reg91 (
      .in(par_done_reg91_in),
      .write_en(par_done_reg91_write_en),
      .clk(clk),
      .out(par_done_reg91_out),
      .done(par_done_reg91_done)
  );
  
  std_reg #(1) par_done_reg92 (
      .in(par_done_reg92_in),
      .write_en(par_done_reg92_write_en),
      .clk(clk),
      .out(par_done_reg92_out),
      .done(par_done_reg92_done)
  );
  
  std_reg #(1) par_done_reg93 (
      .in(par_done_reg93_in),
      .write_en(par_done_reg93_write_en),
      .clk(clk),
      .out(par_done_reg93_out),
      .done(par_done_reg93_done)
  );
  
  std_reg #(1) par_done_reg94 (
      .in(par_done_reg94_in),
      .write_en(par_done_reg94_write_en),
      .clk(clk),
      .out(par_done_reg94_out),
      .done(par_done_reg94_done)
  );
  
  std_reg #(1) par_done_reg95 (
      .in(par_done_reg95_in),
      .write_en(par_done_reg95_write_en),
      .clk(clk),
      .out(par_done_reg95_out),
      .done(par_done_reg95_done)
  );
  
  std_reg #(1) par_done_reg96 (
      .in(par_done_reg96_in),
      .write_en(par_done_reg96_write_en),
      .clk(clk),
      .out(par_done_reg96_out),
      .done(par_done_reg96_done)
  );
  
  std_reg #(1) par_done_reg97 (
      .in(par_done_reg97_in),
      .write_en(par_done_reg97_write_en),
      .clk(clk),
      .out(par_done_reg97_out),
      .done(par_done_reg97_done)
  );
  
  std_reg #(1) par_done_reg98 (
      .in(par_done_reg98_in),
      .write_en(par_done_reg98_write_en),
      .clk(clk),
      .out(par_done_reg98_out),
      .done(par_done_reg98_done)
  );
  
  std_reg #(1) par_done_reg99 (
      .in(par_done_reg99_in),
      .write_en(par_done_reg99_write_en),
      .clk(clk),
      .out(par_done_reg99_out),
      .done(par_done_reg99_done)
  );
  
  std_reg #(1) par_reset10 (
      .in(par_reset10_in),
      .write_en(par_reset10_write_en),
      .clk(clk),
      .out(par_reset10_out),
      .done(par_reset10_done)
  );
  
  std_reg #(1) par_done_reg100 (
      .in(par_done_reg100_in),
      .write_en(par_done_reg100_write_en),
      .clk(clk),
      .out(par_done_reg100_out),
      .done(par_done_reg100_done)
  );
  
  std_reg #(1) par_done_reg101 (
      .in(par_done_reg101_in),
      .write_en(par_done_reg101_write_en),
      .clk(clk),
      .out(par_done_reg101_out),
      .done(par_done_reg101_done)
  );
  
  std_reg #(1) par_done_reg102 (
      .in(par_done_reg102_in),
      .write_en(par_done_reg102_write_en),
      .clk(clk),
      .out(par_done_reg102_out),
      .done(par_done_reg102_done)
  );
  
  std_reg #(1) par_done_reg103 (
      .in(par_done_reg103_in),
      .write_en(par_done_reg103_write_en),
      .clk(clk),
      .out(par_done_reg103_out),
      .done(par_done_reg103_done)
  );
  
  std_reg #(1) par_done_reg104 (
      .in(par_done_reg104_in),
      .write_en(par_done_reg104_write_en),
      .clk(clk),
      .out(par_done_reg104_out),
      .done(par_done_reg104_done)
  );
  
  std_reg #(1) par_done_reg105 (
      .in(par_done_reg105_in),
      .write_en(par_done_reg105_write_en),
      .clk(clk),
      .out(par_done_reg105_out),
      .done(par_done_reg105_done)
  );
  
  std_reg #(1) par_done_reg106 (
      .in(par_done_reg106_in),
      .write_en(par_done_reg106_write_en),
      .clk(clk),
      .out(par_done_reg106_out),
      .done(par_done_reg106_done)
  );
  
  std_reg #(1) par_done_reg107 (
      .in(par_done_reg107_in),
      .write_en(par_done_reg107_write_en),
      .clk(clk),
      .out(par_done_reg107_out),
      .done(par_done_reg107_done)
  );
  
  std_reg #(1) par_done_reg108 (
      .in(par_done_reg108_in),
      .write_en(par_done_reg108_write_en),
      .clk(clk),
      .out(par_done_reg108_out),
      .done(par_done_reg108_done)
  );
  
  std_reg #(1) par_done_reg109 (
      .in(par_done_reg109_in),
      .write_en(par_done_reg109_write_en),
      .clk(clk),
      .out(par_done_reg109_out),
      .done(par_done_reg109_done)
  );
  
  std_reg #(1) par_done_reg110 (
      .in(par_done_reg110_in),
      .write_en(par_done_reg110_write_en),
      .clk(clk),
      .out(par_done_reg110_out),
      .done(par_done_reg110_done)
  );
  
  std_reg #(1) par_done_reg111 (
      .in(par_done_reg111_in),
      .write_en(par_done_reg111_write_en),
      .clk(clk),
      .out(par_done_reg111_out),
      .done(par_done_reg111_done)
  );
  
  std_reg #(1) par_done_reg112 (
      .in(par_done_reg112_in),
      .write_en(par_done_reg112_write_en),
      .clk(clk),
      .out(par_done_reg112_out),
      .done(par_done_reg112_done)
  );
  
  std_reg #(1) par_done_reg113 (
      .in(par_done_reg113_in),
      .write_en(par_done_reg113_write_en),
      .clk(clk),
      .out(par_done_reg113_out),
      .done(par_done_reg113_done)
  );
  
  std_reg #(1) par_done_reg114 (
      .in(par_done_reg114_in),
      .write_en(par_done_reg114_write_en),
      .clk(clk),
      .out(par_done_reg114_out),
      .done(par_done_reg114_done)
  );
  
  std_reg #(1) par_done_reg115 (
      .in(par_done_reg115_in),
      .write_en(par_done_reg115_write_en),
      .clk(clk),
      .out(par_done_reg115_out),
      .done(par_done_reg115_done)
  );
  
  std_reg #(1) par_done_reg116 (
      .in(par_done_reg116_in),
      .write_en(par_done_reg116_write_en),
      .clk(clk),
      .out(par_done_reg116_out),
      .done(par_done_reg116_done)
  );
  
  std_reg #(1) par_done_reg117 (
      .in(par_done_reg117_in),
      .write_en(par_done_reg117_write_en),
      .clk(clk),
      .out(par_done_reg117_out),
      .done(par_done_reg117_done)
  );
  
  std_reg #(1) par_done_reg118 (
      .in(par_done_reg118_in),
      .write_en(par_done_reg118_write_en),
      .clk(clk),
      .out(par_done_reg118_out),
      .done(par_done_reg118_done)
  );
  
  std_reg #(1) par_done_reg119 (
      .in(par_done_reg119_in),
      .write_en(par_done_reg119_write_en),
      .clk(clk),
      .out(par_done_reg119_out),
      .done(par_done_reg119_done)
  );
  
  std_reg #(1) par_done_reg120 (
      .in(par_done_reg120_in),
      .write_en(par_done_reg120_write_en),
      .clk(clk),
      .out(par_done_reg120_out),
      .done(par_done_reg120_done)
  );
  
  std_reg #(1) par_done_reg121 (
      .in(par_done_reg121_in),
      .write_en(par_done_reg121_write_en),
      .clk(clk),
      .out(par_done_reg121_out),
      .done(par_done_reg121_done)
  );
  
  std_reg #(1) par_done_reg122 (
      .in(par_done_reg122_in),
      .write_en(par_done_reg122_write_en),
      .clk(clk),
      .out(par_done_reg122_out),
      .done(par_done_reg122_done)
  );
  
  std_reg #(1) par_done_reg123 (
      .in(par_done_reg123_in),
      .write_en(par_done_reg123_write_en),
      .clk(clk),
      .out(par_done_reg123_out),
      .done(par_done_reg123_done)
  );
  
  std_reg #(1) par_done_reg124 (
      .in(par_done_reg124_in),
      .write_en(par_done_reg124_write_en),
      .clk(clk),
      .out(par_done_reg124_out),
      .done(par_done_reg124_done)
  );
  
  std_reg #(1) par_done_reg125 (
      .in(par_done_reg125_in),
      .write_en(par_done_reg125_write_en),
      .clk(clk),
      .out(par_done_reg125_out),
      .done(par_done_reg125_done)
  );
  
  std_reg #(1) par_done_reg126 (
      .in(par_done_reg126_in),
      .write_en(par_done_reg126_write_en),
      .clk(clk),
      .out(par_done_reg126_out),
      .done(par_done_reg126_done)
  );
  
  std_reg #(1) par_done_reg127 (
      .in(par_done_reg127_in),
      .write_en(par_done_reg127_write_en),
      .clk(clk),
      .out(par_done_reg127_out),
      .done(par_done_reg127_done)
  );
  
  std_reg #(1) par_done_reg128 (
      .in(par_done_reg128_in),
      .write_en(par_done_reg128_write_en),
      .clk(clk),
      .out(par_done_reg128_out),
      .done(par_done_reg128_done)
  );
  
  std_reg #(1) par_done_reg129 (
      .in(par_done_reg129_in),
      .write_en(par_done_reg129_write_en),
      .clk(clk),
      .out(par_done_reg129_out),
      .done(par_done_reg129_done)
  );
  
  std_reg #(1) par_reset11 (
      .in(par_reset11_in),
      .write_en(par_reset11_write_en),
      .clk(clk),
      .out(par_reset11_out),
      .done(par_reset11_done)
  );
  
  std_reg #(1) par_done_reg130 (
      .in(par_done_reg130_in),
      .write_en(par_done_reg130_write_en),
      .clk(clk),
      .out(par_done_reg130_out),
      .done(par_done_reg130_done)
  );
  
  std_reg #(1) par_done_reg131 (
      .in(par_done_reg131_in),
      .write_en(par_done_reg131_write_en),
      .clk(clk),
      .out(par_done_reg131_out),
      .done(par_done_reg131_done)
  );
  
  std_reg #(1) par_done_reg132 (
      .in(par_done_reg132_in),
      .write_en(par_done_reg132_write_en),
      .clk(clk),
      .out(par_done_reg132_out),
      .done(par_done_reg132_done)
  );
  
  std_reg #(1) par_done_reg133 (
      .in(par_done_reg133_in),
      .write_en(par_done_reg133_write_en),
      .clk(clk),
      .out(par_done_reg133_out),
      .done(par_done_reg133_done)
  );
  
  std_reg #(1) par_done_reg134 (
      .in(par_done_reg134_in),
      .write_en(par_done_reg134_write_en),
      .clk(clk),
      .out(par_done_reg134_out),
      .done(par_done_reg134_done)
  );
  
  std_reg #(1) par_done_reg135 (
      .in(par_done_reg135_in),
      .write_en(par_done_reg135_write_en),
      .clk(clk),
      .out(par_done_reg135_out),
      .done(par_done_reg135_done)
  );
  
  std_reg #(1) par_done_reg136 (
      .in(par_done_reg136_in),
      .write_en(par_done_reg136_write_en),
      .clk(clk),
      .out(par_done_reg136_out),
      .done(par_done_reg136_done)
  );
  
  std_reg #(1) par_done_reg137 (
      .in(par_done_reg137_in),
      .write_en(par_done_reg137_write_en),
      .clk(clk),
      .out(par_done_reg137_out),
      .done(par_done_reg137_done)
  );
  
  std_reg #(1) par_done_reg138 (
      .in(par_done_reg138_in),
      .write_en(par_done_reg138_write_en),
      .clk(clk),
      .out(par_done_reg138_out),
      .done(par_done_reg138_done)
  );
  
  std_reg #(1) par_done_reg139 (
      .in(par_done_reg139_in),
      .write_en(par_done_reg139_write_en),
      .clk(clk),
      .out(par_done_reg139_out),
      .done(par_done_reg139_done)
  );
  
  std_reg #(1) par_done_reg140 (
      .in(par_done_reg140_in),
      .write_en(par_done_reg140_write_en),
      .clk(clk),
      .out(par_done_reg140_out),
      .done(par_done_reg140_done)
  );
  
  std_reg #(1) par_done_reg141 (
      .in(par_done_reg141_in),
      .write_en(par_done_reg141_write_en),
      .clk(clk),
      .out(par_done_reg141_out),
      .done(par_done_reg141_done)
  );
  
  std_reg #(1) par_done_reg142 (
      .in(par_done_reg142_in),
      .write_en(par_done_reg142_write_en),
      .clk(clk),
      .out(par_done_reg142_out),
      .done(par_done_reg142_done)
  );
  
  std_reg #(1) par_done_reg143 (
      .in(par_done_reg143_in),
      .write_en(par_done_reg143_write_en),
      .clk(clk),
      .out(par_done_reg143_out),
      .done(par_done_reg143_done)
  );
  
  std_reg #(1) par_done_reg144 (
      .in(par_done_reg144_in),
      .write_en(par_done_reg144_write_en),
      .clk(clk),
      .out(par_done_reg144_out),
      .done(par_done_reg144_done)
  );
  
  std_reg #(1) par_done_reg145 (
      .in(par_done_reg145_in),
      .write_en(par_done_reg145_write_en),
      .clk(clk),
      .out(par_done_reg145_out),
      .done(par_done_reg145_done)
  );
  
  std_reg #(1) par_done_reg146 (
      .in(par_done_reg146_in),
      .write_en(par_done_reg146_write_en),
      .clk(clk),
      .out(par_done_reg146_out),
      .done(par_done_reg146_done)
  );
  
  std_reg #(1) par_done_reg147 (
      .in(par_done_reg147_in),
      .write_en(par_done_reg147_write_en),
      .clk(clk),
      .out(par_done_reg147_out),
      .done(par_done_reg147_done)
  );
  
  std_reg #(1) par_done_reg148 (
      .in(par_done_reg148_in),
      .write_en(par_done_reg148_write_en),
      .clk(clk),
      .out(par_done_reg148_out),
      .done(par_done_reg148_done)
  );
  
  std_reg #(1) par_done_reg149 (
      .in(par_done_reg149_in),
      .write_en(par_done_reg149_write_en),
      .clk(clk),
      .out(par_done_reg149_out),
      .done(par_done_reg149_done)
  );
  
  std_reg #(1) par_done_reg150 (
      .in(par_done_reg150_in),
      .write_en(par_done_reg150_write_en),
      .clk(clk),
      .out(par_done_reg150_out),
      .done(par_done_reg150_done)
  );
  
  std_reg #(1) par_done_reg151 (
      .in(par_done_reg151_in),
      .write_en(par_done_reg151_write_en),
      .clk(clk),
      .out(par_done_reg151_out),
      .done(par_done_reg151_done)
  );
  
  std_reg #(1) par_done_reg152 (
      .in(par_done_reg152_in),
      .write_en(par_done_reg152_write_en),
      .clk(clk),
      .out(par_done_reg152_out),
      .done(par_done_reg152_done)
  );
  
  std_reg #(1) par_reset12 (
      .in(par_reset12_in),
      .write_en(par_reset12_write_en),
      .clk(clk),
      .out(par_reset12_out),
      .done(par_reset12_done)
  );
  
  std_reg #(1) par_done_reg153 (
      .in(par_done_reg153_in),
      .write_en(par_done_reg153_write_en),
      .clk(clk),
      .out(par_done_reg153_out),
      .done(par_done_reg153_done)
  );
  
  std_reg #(1) par_done_reg154 (
      .in(par_done_reg154_in),
      .write_en(par_done_reg154_write_en),
      .clk(clk),
      .out(par_done_reg154_out),
      .done(par_done_reg154_done)
  );
  
  std_reg #(1) par_done_reg155 (
      .in(par_done_reg155_in),
      .write_en(par_done_reg155_write_en),
      .clk(clk),
      .out(par_done_reg155_out),
      .done(par_done_reg155_done)
  );
  
  std_reg #(1) par_done_reg156 (
      .in(par_done_reg156_in),
      .write_en(par_done_reg156_write_en),
      .clk(clk),
      .out(par_done_reg156_out),
      .done(par_done_reg156_done)
  );
  
  std_reg #(1) par_done_reg157 (
      .in(par_done_reg157_in),
      .write_en(par_done_reg157_write_en),
      .clk(clk),
      .out(par_done_reg157_out),
      .done(par_done_reg157_done)
  );
  
  std_reg #(1) par_done_reg158 (
      .in(par_done_reg158_in),
      .write_en(par_done_reg158_write_en),
      .clk(clk),
      .out(par_done_reg158_out),
      .done(par_done_reg158_done)
  );
  
  std_reg #(1) par_done_reg159 (
      .in(par_done_reg159_in),
      .write_en(par_done_reg159_write_en),
      .clk(clk),
      .out(par_done_reg159_out),
      .done(par_done_reg159_done)
  );
  
  std_reg #(1) par_done_reg160 (
      .in(par_done_reg160_in),
      .write_en(par_done_reg160_write_en),
      .clk(clk),
      .out(par_done_reg160_out),
      .done(par_done_reg160_done)
  );
  
  std_reg #(1) par_done_reg161 (
      .in(par_done_reg161_in),
      .write_en(par_done_reg161_write_en),
      .clk(clk),
      .out(par_done_reg161_out),
      .done(par_done_reg161_done)
  );
  
  std_reg #(1) par_done_reg162 (
      .in(par_done_reg162_in),
      .write_en(par_done_reg162_write_en),
      .clk(clk),
      .out(par_done_reg162_out),
      .done(par_done_reg162_done)
  );
  
  std_reg #(1) par_done_reg163 (
      .in(par_done_reg163_in),
      .write_en(par_done_reg163_write_en),
      .clk(clk),
      .out(par_done_reg163_out),
      .done(par_done_reg163_done)
  );
  
  std_reg #(1) par_done_reg164 (
      .in(par_done_reg164_in),
      .write_en(par_done_reg164_write_en),
      .clk(clk),
      .out(par_done_reg164_out),
      .done(par_done_reg164_done)
  );
  
  std_reg #(1) par_done_reg165 (
      .in(par_done_reg165_in),
      .write_en(par_done_reg165_write_en),
      .clk(clk),
      .out(par_done_reg165_out),
      .done(par_done_reg165_done)
  );
  
  std_reg #(1) par_done_reg166 (
      .in(par_done_reg166_in),
      .write_en(par_done_reg166_write_en),
      .clk(clk),
      .out(par_done_reg166_out),
      .done(par_done_reg166_done)
  );
  
  std_reg #(1) par_done_reg167 (
      .in(par_done_reg167_in),
      .write_en(par_done_reg167_write_en),
      .clk(clk),
      .out(par_done_reg167_out),
      .done(par_done_reg167_done)
  );
  
  std_reg #(1) par_done_reg168 (
      .in(par_done_reg168_in),
      .write_en(par_done_reg168_write_en),
      .clk(clk),
      .out(par_done_reg168_out),
      .done(par_done_reg168_done)
  );
  
  std_reg #(1) par_done_reg169 (
      .in(par_done_reg169_in),
      .write_en(par_done_reg169_write_en),
      .clk(clk),
      .out(par_done_reg169_out),
      .done(par_done_reg169_done)
  );
  
  std_reg #(1) par_done_reg170 (
      .in(par_done_reg170_in),
      .write_en(par_done_reg170_write_en),
      .clk(clk),
      .out(par_done_reg170_out),
      .done(par_done_reg170_done)
  );
  
  std_reg #(1) par_done_reg171 (
      .in(par_done_reg171_in),
      .write_en(par_done_reg171_write_en),
      .clk(clk),
      .out(par_done_reg171_out),
      .done(par_done_reg171_done)
  );
  
  std_reg #(1) par_done_reg172 (
      .in(par_done_reg172_in),
      .write_en(par_done_reg172_write_en),
      .clk(clk),
      .out(par_done_reg172_out),
      .done(par_done_reg172_done)
  );
  
  std_reg #(1) par_done_reg173 (
      .in(par_done_reg173_in),
      .write_en(par_done_reg173_write_en),
      .clk(clk),
      .out(par_done_reg173_out),
      .done(par_done_reg173_done)
  );
  
  std_reg #(1) par_done_reg174 (
      .in(par_done_reg174_in),
      .write_en(par_done_reg174_write_en),
      .clk(clk),
      .out(par_done_reg174_out),
      .done(par_done_reg174_done)
  );
  
  std_reg #(1) par_done_reg175 (
      .in(par_done_reg175_in),
      .write_en(par_done_reg175_write_en),
      .clk(clk),
      .out(par_done_reg175_out),
      .done(par_done_reg175_done)
  );
  
  std_reg #(1) par_done_reg176 (
      .in(par_done_reg176_in),
      .write_en(par_done_reg176_write_en),
      .clk(clk),
      .out(par_done_reg176_out),
      .done(par_done_reg176_done)
  );
  
  std_reg #(1) par_done_reg177 (
      .in(par_done_reg177_in),
      .write_en(par_done_reg177_write_en),
      .clk(clk),
      .out(par_done_reg177_out),
      .done(par_done_reg177_done)
  );
  
  std_reg #(1) par_done_reg178 (
      .in(par_done_reg178_in),
      .write_en(par_done_reg178_write_en),
      .clk(clk),
      .out(par_done_reg178_out),
      .done(par_done_reg178_done)
  );
  
  std_reg #(1) par_done_reg179 (
      .in(par_done_reg179_in),
      .write_en(par_done_reg179_write_en),
      .clk(clk),
      .out(par_done_reg179_out),
      .done(par_done_reg179_done)
  );
  
  std_reg #(1) par_done_reg180 (
      .in(par_done_reg180_in),
      .write_en(par_done_reg180_write_en),
      .clk(clk),
      .out(par_done_reg180_out),
      .done(par_done_reg180_done)
  );
  
  std_reg #(1) par_done_reg181 (
      .in(par_done_reg181_in),
      .write_en(par_done_reg181_write_en),
      .clk(clk),
      .out(par_done_reg181_out),
      .done(par_done_reg181_done)
  );
  
  std_reg #(1) par_done_reg182 (
      .in(par_done_reg182_in),
      .write_en(par_done_reg182_write_en),
      .clk(clk),
      .out(par_done_reg182_out),
      .done(par_done_reg182_done)
  );
  
  std_reg #(1) par_done_reg183 (
      .in(par_done_reg183_in),
      .write_en(par_done_reg183_write_en),
      .clk(clk),
      .out(par_done_reg183_out),
      .done(par_done_reg183_done)
  );
  
  std_reg #(1) par_done_reg184 (
      .in(par_done_reg184_in),
      .write_en(par_done_reg184_write_en),
      .clk(clk),
      .out(par_done_reg184_out),
      .done(par_done_reg184_done)
  );
  
  std_reg #(1) par_done_reg185 (
      .in(par_done_reg185_in),
      .write_en(par_done_reg185_write_en),
      .clk(clk),
      .out(par_done_reg185_out),
      .done(par_done_reg185_done)
  );
  
  std_reg #(1) par_done_reg186 (
      .in(par_done_reg186_in),
      .write_en(par_done_reg186_write_en),
      .clk(clk),
      .out(par_done_reg186_out),
      .done(par_done_reg186_done)
  );
  
  std_reg #(1) par_done_reg187 (
      .in(par_done_reg187_in),
      .write_en(par_done_reg187_write_en),
      .clk(clk),
      .out(par_done_reg187_out),
      .done(par_done_reg187_done)
  );
  
  std_reg #(1) par_done_reg188 (
      .in(par_done_reg188_in),
      .write_en(par_done_reg188_write_en),
      .clk(clk),
      .out(par_done_reg188_out),
      .done(par_done_reg188_done)
  );
  
  std_reg #(1) par_reset13 (
      .in(par_reset13_in),
      .write_en(par_reset13_write_en),
      .clk(clk),
      .out(par_reset13_out),
      .done(par_reset13_done)
  );
  
  std_reg #(1) par_done_reg189 (
      .in(par_done_reg189_in),
      .write_en(par_done_reg189_write_en),
      .clk(clk),
      .out(par_done_reg189_out),
      .done(par_done_reg189_done)
  );
  
  std_reg #(1) par_done_reg190 (
      .in(par_done_reg190_in),
      .write_en(par_done_reg190_write_en),
      .clk(clk),
      .out(par_done_reg190_out),
      .done(par_done_reg190_done)
  );
  
  std_reg #(1) par_done_reg191 (
      .in(par_done_reg191_in),
      .write_en(par_done_reg191_write_en),
      .clk(clk),
      .out(par_done_reg191_out),
      .done(par_done_reg191_done)
  );
  
  std_reg #(1) par_done_reg192 (
      .in(par_done_reg192_in),
      .write_en(par_done_reg192_write_en),
      .clk(clk),
      .out(par_done_reg192_out),
      .done(par_done_reg192_done)
  );
  
  std_reg #(1) par_done_reg193 (
      .in(par_done_reg193_in),
      .write_en(par_done_reg193_write_en),
      .clk(clk),
      .out(par_done_reg193_out),
      .done(par_done_reg193_done)
  );
  
  std_reg #(1) par_done_reg194 (
      .in(par_done_reg194_in),
      .write_en(par_done_reg194_write_en),
      .clk(clk),
      .out(par_done_reg194_out),
      .done(par_done_reg194_done)
  );
  
  std_reg #(1) par_done_reg195 (
      .in(par_done_reg195_in),
      .write_en(par_done_reg195_write_en),
      .clk(clk),
      .out(par_done_reg195_out),
      .done(par_done_reg195_done)
  );
  
  std_reg #(1) par_done_reg196 (
      .in(par_done_reg196_in),
      .write_en(par_done_reg196_write_en),
      .clk(clk),
      .out(par_done_reg196_out),
      .done(par_done_reg196_done)
  );
  
  std_reg #(1) par_done_reg197 (
      .in(par_done_reg197_in),
      .write_en(par_done_reg197_write_en),
      .clk(clk),
      .out(par_done_reg197_out),
      .done(par_done_reg197_done)
  );
  
  std_reg #(1) par_done_reg198 (
      .in(par_done_reg198_in),
      .write_en(par_done_reg198_write_en),
      .clk(clk),
      .out(par_done_reg198_out),
      .done(par_done_reg198_done)
  );
  
  std_reg #(1) par_done_reg199 (
      .in(par_done_reg199_in),
      .write_en(par_done_reg199_write_en),
      .clk(clk),
      .out(par_done_reg199_out),
      .done(par_done_reg199_done)
  );
  
  std_reg #(1) par_done_reg200 (
      .in(par_done_reg200_in),
      .write_en(par_done_reg200_write_en),
      .clk(clk),
      .out(par_done_reg200_out),
      .done(par_done_reg200_done)
  );
  
  std_reg #(1) par_done_reg201 (
      .in(par_done_reg201_in),
      .write_en(par_done_reg201_write_en),
      .clk(clk),
      .out(par_done_reg201_out),
      .done(par_done_reg201_done)
  );
  
  std_reg #(1) par_done_reg202 (
      .in(par_done_reg202_in),
      .write_en(par_done_reg202_write_en),
      .clk(clk),
      .out(par_done_reg202_out),
      .done(par_done_reg202_done)
  );
  
  std_reg #(1) par_done_reg203 (
      .in(par_done_reg203_in),
      .write_en(par_done_reg203_write_en),
      .clk(clk),
      .out(par_done_reg203_out),
      .done(par_done_reg203_done)
  );
  
  std_reg #(1) par_done_reg204 (
      .in(par_done_reg204_in),
      .write_en(par_done_reg204_write_en),
      .clk(clk),
      .out(par_done_reg204_out),
      .done(par_done_reg204_done)
  );
  
  std_reg #(1) par_done_reg205 (
      .in(par_done_reg205_in),
      .write_en(par_done_reg205_write_en),
      .clk(clk),
      .out(par_done_reg205_out),
      .done(par_done_reg205_done)
  );
  
  std_reg #(1) par_done_reg206 (
      .in(par_done_reg206_in),
      .write_en(par_done_reg206_write_en),
      .clk(clk),
      .out(par_done_reg206_out),
      .done(par_done_reg206_done)
  );
  
  std_reg #(1) par_done_reg207 (
      .in(par_done_reg207_in),
      .write_en(par_done_reg207_write_en),
      .clk(clk),
      .out(par_done_reg207_out),
      .done(par_done_reg207_done)
  );
  
  std_reg #(1) par_done_reg208 (
      .in(par_done_reg208_in),
      .write_en(par_done_reg208_write_en),
      .clk(clk),
      .out(par_done_reg208_out),
      .done(par_done_reg208_done)
  );
  
  std_reg #(1) par_done_reg209 (
      .in(par_done_reg209_in),
      .write_en(par_done_reg209_write_en),
      .clk(clk),
      .out(par_done_reg209_out),
      .done(par_done_reg209_done)
  );
  
  std_reg #(1) par_done_reg210 (
      .in(par_done_reg210_in),
      .write_en(par_done_reg210_write_en),
      .clk(clk),
      .out(par_done_reg210_out),
      .done(par_done_reg210_done)
  );
  
  std_reg #(1) par_done_reg211 (
      .in(par_done_reg211_in),
      .write_en(par_done_reg211_write_en),
      .clk(clk),
      .out(par_done_reg211_out),
      .done(par_done_reg211_done)
  );
  
  std_reg #(1) par_done_reg212 (
      .in(par_done_reg212_in),
      .write_en(par_done_reg212_write_en),
      .clk(clk),
      .out(par_done_reg212_out),
      .done(par_done_reg212_done)
  );
  
  std_reg #(1) par_reset14 (
      .in(par_reset14_in),
      .write_en(par_reset14_write_en),
      .clk(clk),
      .out(par_reset14_out),
      .done(par_reset14_done)
  );
  
  std_reg #(1) par_done_reg213 (
      .in(par_done_reg213_in),
      .write_en(par_done_reg213_write_en),
      .clk(clk),
      .out(par_done_reg213_out),
      .done(par_done_reg213_done)
  );
  
  std_reg #(1) par_done_reg214 (
      .in(par_done_reg214_in),
      .write_en(par_done_reg214_write_en),
      .clk(clk),
      .out(par_done_reg214_out),
      .done(par_done_reg214_done)
  );
  
  std_reg #(1) par_done_reg215 (
      .in(par_done_reg215_in),
      .write_en(par_done_reg215_write_en),
      .clk(clk),
      .out(par_done_reg215_out),
      .done(par_done_reg215_done)
  );
  
  std_reg #(1) par_done_reg216 (
      .in(par_done_reg216_in),
      .write_en(par_done_reg216_write_en),
      .clk(clk),
      .out(par_done_reg216_out),
      .done(par_done_reg216_done)
  );
  
  std_reg #(1) par_done_reg217 (
      .in(par_done_reg217_in),
      .write_en(par_done_reg217_write_en),
      .clk(clk),
      .out(par_done_reg217_out),
      .done(par_done_reg217_done)
  );
  
  std_reg #(1) par_done_reg218 (
      .in(par_done_reg218_in),
      .write_en(par_done_reg218_write_en),
      .clk(clk),
      .out(par_done_reg218_out),
      .done(par_done_reg218_done)
  );
  
  std_reg #(1) par_done_reg219 (
      .in(par_done_reg219_in),
      .write_en(par_done_reg219_write_en),
      .clk(clk),
      .out(par_done_reg219_out),
      .done(par_done_reg219_done)
  );
  
  std_reg #(1) par_done_reg220 (
      .in(par_done_reg220_in),
      .write_en(par_done_reg220_write_en),
      .clk(clk),
      .out(par_done_reg220_out),
      .done(par_done_reg220_done)
  );
  
  std_reg #(1) par_done_reg221 (
      .in(par_done_reg221_in),
      .write_en(par_done_reg221_write_en),
      .clk(clk),
      .out(par_done_reg221_out),
      .done(par_done_reg221_done)
  );
  
  std_reg #(1) par_done_reg222 (
      .in(par_done_reg222_in),
      .write_en(par_done_reg222_write_en),
      .clk(clk),
      .out(par_done_reg222_out),
      .done(par_done_reg222_done)
  );
  
  std_reg #(1) par_done_reg223 (
      .in(par_done_reg223_in),
      .write_en(par_done_reg223_write_en),
      .clk(clk),
      .out(par_done_reg223_out),
      .done(par_done_reg223_done)
  );
  
  std_reg #(1) par_done_reg224 (
      .in(par_done_reg224_in),
      .write_en(par_done_reg224_write_en),
      .clk(clk),
      .out(par_done_reg224_out),
      .done(par_done_reg224_done)
  );
  
  std_reg #(1) par_done_reg225 (
      .in(par_done_reg225_in),
      .write_en(par_done_reg225_write_en),
      .clk(clk),
      .out(par_done_reg225_out),
      .done(par_done_reg225_done)
  );
  
  std_reg #(1) par_done_reg226 (
      .in(par_done_reg226_in),
      .write_en(par_done_reg226_write_en),
      .clk(clk),
      .out(par_done_reg226_out),
      .done(par_done_reg226_done)
  );
  
  std_reg #(1) par_done_reg227 (
      .in(par_done_reg227_in),
      .write_en(par_done_reg227_write_en),
      .clk(clk),
      .out(par_done_reg227_out),
      .done(par_done_reg227_done)
  );
  
  std_reg #(1) par_done_reg228 (
      .in(par_done_reg228_in),
      .write_en(par_done_reg228_write_en),
      .clk(clk),
      .out(par_done_reg228_out),
      .done(par_done_reg228_done)
  );
  
  std_reg #(1) par_done_reg229 (
      .in(par_done_reg229_in),
      .write_en(par_done_reg229_write_en),
      .clk(clk),
      .out(par_done_reg229_out),
      .done(par_done_reg229_done)
  );
  
  std_reg #(1) par_done_reg230 (
      .in(par_done_reg230_in),
      .write_en(par_done_reg230_write_en),
      .clk(clk),
      .out(par_done_reg230_out),
      .done(par_done_reg230_done)
  );
  
  std_reg #(1) par_done_reg231 (
      .in(par_done_reg231_in),
      .write_en(par_done_reg231_write_en),
      .clk(clk),
      .out(par_done_reg231_out),
      .done(par_done_reg231_done)
  );
  
  std_reg #(1) par_done_reg232 (
      .in(par_done_reg232_in),
      .write_en(par_done_reg232_write_en),
      .clk(clk),
      .out(par_done_reg232_out),
      .done(par_done_reg232_done)
  );
  
  std_reg #(1) par_done_reg233 (
      .in(par_done_reg233_in),
      .write_en(par_done_reg233_write_en),
      .clk(clk),
      .out(par_done_reg233_out),
      .done(par_done_reg233_done)
  );
  
  std_reg #(1) par_done_reg234 (
      .in(par_done_reg234_in),
      .write_en(par_done_reg234_write_en),
      .clk(clk),
      .out(par_done_reg234_out),
      .done(par_done_reg234_done)
  );
  
  std_reg #(1) par_done_reg235 (
      .in(par_done_reg235_in),
      .write_en(par_done_reg235_write_en),
      .clk(clk),
      .out(par_done_reg235_out),
      .done(par_done_reg235_done)
  );
  
  std_reg #(1) par_done_reg236 (
      .in(par_done_reg236_in),
      .write_en(par_done_reg236_write_en),
      .clk(clk),
      .out(par_done_reg236_out),
      .done(par_done_reg236_done)
  );
  
  std_reg #(1) par_done_reg237 (
      .in(par_done_reg237_in),
      .write_en(par_done_reg237_write_en),
      .clk(clk),
      .out(par_done_reg237_out),
      .done(par_done_reg237_done)
  );
  
  std_reg #(1) par_done_reg238 (
      .in(par_done_reg238_in),
      .write_en(par_done_reg238_write_en),
      .clk(clk),
      .out(par_done_reg238_out),
      .done(par_done_reg238_done)
  );
  
  std_reg #(1) par_done_reg239 (
      .in(par_done_reg239_in),
      .write_en(par_done_reg239_write_en),
      .clk(clk),
      .out(par_done_reg239_out),
      .done(par_done_reg239_done)
  );
  
  std_reg #(1) par_done_reg240 (
      .in(par_done_reg240_in),
      .write_en(par_done_reg240_write_en),
      .clk(clk),
      .out(par_done_reg240_out),
      .done(par_done_reg240_done)
  );
  
  std_reg #(1) par_done_reg241 (
      .in(par_done_reg241_in),
      .write_en(par_done_reg241_write_en),
      .clk(clk),
      .out(par_done_reg241_out),
      .done(par_done_reg241_done)
  );
  
  std_reg #(1) par_done_reg242 (
      .in(par_done_reg242_in),
      .write_en(par_done_reg242_write_en),
      .clk(clk),
      .out(par_done_reg242_out),
      .done(par_done_reg242_done)
  );
  
  std_reg #(1) par_done_reg243 (
      .in(par_done_reg243_in),
      .write_en(par_done_reg243_write_en),
      .clk(clk),
      .out(par_done_reg243_out),
      .done(par_done_reg243_done)
  );
  
  std_reg #(1) par_done_reg244 (
      .in(par_done_reg244_in),
      .write_en(par_done_reg244_write_en),
      .clk(clk),
      .out(par_done_reg244_out),
      .done(par_done_reg244_done)
  );
  
  std_reg #(1) par_done_reg245 (
      .in(par_done_reg245_in),
      .write_en(par_done_reg245_write_en),
      .clk(clk),
      .out(par_done_reg245_out),
      .done(par_done_reg245_done)
  );
  
  std_reg #(1) par_done_reg246 (
      .in(par_done_reg246_in),
      .write_en(par_done_reg246_write_en),
      .clk(clk),
      .out(par_done_reg246_out),
      .done(par_done_reg246_done)
  );
  
  std_reg #(1) par_done_reg247 (
      .in(par_done_reg247_in),
      .write_en(par_done_reg247_write_en),
      .clk(clk),
      .out(par_done_reg247_out),
      .done(par_done_reg247_done)
  );
  
  std_reg #(1) par_done_reg248 (
      .in(par_done_reg248_in),
      .write_en(par_done_reg248_write_en),
      .clk(clk),
      .out(par_done_reg248_out),
      .done(par_done_reg248_done)
  );
  
  std_reg #(1) par_done_reg249 (
      .in(par_done_reg249_in),
      .write_en(par_done_reg249_write_en),
      .clk(clk),
      .out(par_done_reg249_out),
      .done(par_done_reg249_done)
  );
  
  std_reg #(1) par_done_reg250 (
      .in(par_done_reg250_in),
      .write_en(par_done_reg250_write_en),
      .clk(clk),
      .out(par_done_reg250_out),
      .done(par_done_reg250_done)
  );
  
  std_reg #(1) par_reset15 (
      .in(par_reset15_in),
      .write_en(par_reset15_write_en),
      .clk(clk),
      .out(par_reset15_out),
      .done(par_reset15_done)
  );
  
  std_reg #(1) par_done_reg251 (
      .in(par_done_reg251_in),
      .write_en(par_done_reg251_write_en),
      .clk(clk),
      .out(par_done_reg251_out),
      .done(par_done_reg251_done)
  );
  
  std_reg #(1) par_done_reg252 (
      .in(par_done_reg252_in),
      .write_en(par_done_reg252_write_en),
      .clk(clk),
      .out(par_done_reg252_out),
      .done(par_done_reg252_done)
  );
  
  std_reg #(1) par_done_reg253 (
      .in(par_done_reg253_in),
      .write_en(par_done_reg253_write_en),
      .clk(clk),
      .out(par_done_reg253_out),
      .done(par_done_reg253_done)
  );
  
  std_reg #(1) par_done_reg254 (
      .in(par_done_reg254_in),
      .write_en(par_done_reg254_write_en),
      .clk(clk),
      .out(par_done_reg254_out),
      .done(par_done_reg254_done)
  );
  
  std_reg #(1) par_done_reg255 (
      .in(par_done_reg255_in),
      .write_en(par_done_reg255_write_en),
      .clk(clk),
      .out(par_done_reg255_out),
      .done(par_done_reg255_done)
  );
  
  std_reg #(1) par_done_reg256 (
      .in(par_done_reg256_in),
      .write_en(par_done_reg256_write_en),
      .clk(clk),
      .out(par_done_reg256_out),
      .done(par_done_reg256_done)
  );
  
  std_reg #(1) par_done_reg257 (
      .in(par_done_reg257_in),
      .write_en(par_done_reg257_write_en),
      .clk(clk),
      .out(par_done_reg257_out),
      .done(par_done_reg257_done)
  );
  
  std_reg #(1) par_done_reg258 (
      .in(par_done_reg258_in),
      .write_en(par_done_reg258_write_en),
      .clk(clk),
      .out(par_done_reg258_out),
      .done(par_done_reg258_done)
  );
  
  std_reg #(1) par_done_reg259 (
      .in(par_done_reg259_in),
      .write_en(par_done_reg259_write_en),
      .clk(clk),
      .out(par_done_reg259_out),
      .done(par_done_reg259_done)
  );
  
  std_reg #(1) par_done_reg260 (
      .in(par_done_reg260_in),
      .write_en(par_done_reg260_write_en),
      .clk(clk),
      .out(par_done_reg260_out),
      .done(par_done_reg260_done)
  );
  
  std_reg #(1) par_done_reg261 (
      .in(par_done_reg261_in),
      .write_en(par_done_reg261_write_en),
      .clk(clk),
      .out(par_done_reg261_out),
      .done(par_done_reg261_done)
  );
  
  std_reg #(1) par_done_reg262 (
      .in(par_done_reg262_in),
      .write_en(par_done_reg262_write_en),
      .clk(clk),
      .out(par_done_reg262_out),
      .done(par_done_reg262_done)
  );
  
  std_reg #(1) par_done_reg263 (
      .in(par_done_reg263_in),
      .write_en(par_done_reg263_write_en),
      .clk(clk),
      .out(par_done_reg263_out),
      .done(par_done_reg263_done)
  );
  
  std_reg #(1) par_done_reg264 (
      .in(par_done_reg264_in),
      .write_en(par_done_reg264_write_en),
      .clk(clk),
      .out(par_done_reg264_out),
      .done(par_done_reg264_done)
  );
  
  std_reg #(1) par_done_reg265 (
      .in(par_done_reg265_in),
      .write_en(par_done_reg265_write_en),
      .clk(clk),
      .out(par_done_reg265_out),
      .done(par_done_reg265_done)
  );
  
  std_reg #(1) par_done_reg266 (
      .in(par_done_reg266_in),
      .write_en(par_done_reg266_write_en),
      .clk(clk),
      .out(par_done_reg266_out),
      .done(par_done_reg266_done)
  );
  
  std_reg #(1) par_done_reg267 (
      .in(par_done_reg267_in),
      .write_en(par_done_reg267_write_en),
      .clk(clk),
      .out(par_done_reg267_out),
      .done(par_done_reg267_done)
  );
  
  std_reg #(1) par_done_reg268 (
      .in(par_done_reg268_in),
      .write_en(par_done_reg268_write_en),
      .clk(clk),
      .out(par_done_reg268_out),
      .done(par_done_reg268_done)
  );
  
  std_reg #(1) par_done_reg269 (
      .in(par_done_reg269_in),
      .write_en(par_done_reg269_write_en),
      .clk(clk),
      .out(par_done_reg269_out),
      .done(par_done_reg269_done)
  );
  
  std_reg #(1) par_done_reg270 (
      .in(par_done_reg270_in),
      .write_en(par_done_reg270_write_en),
      .clk(clk),
      .out(par_done_reg270_out),
      .done(par_done_reg270_done)
  );
  
  std_reg #(1) par_done_reg271 (
      .in(par_done_reg271_in),
      .write_en(par_done_reg271_write_en),
      .clk(clk),
      .out(par_done_reg271_out),
      .done(par_done_reg271_done)
  );
  
  std_reg #(1) par_done_reg272 (
      .in(par_done_reg272_in),
      .write_en(par_done_reg272_write_en),
      .clk(clk),
      .out(par_done_reg272_out),
      .done(par_done_reg272_done)
  );
  
  std_reg #(1) par_done_reg273 (
      .in(par_done_reg273_in),
      .write_en(par_done_reg273_write_en),
      .clk(clk),
      .out(par_done_reg273_out),
      .done(par_done_reg273_done)
  );
  
  std_reg #(1) par_reset16 (
      .in(par_reset16_in),
      .write_en(par_reset16_write_en),
      .clk(clk),
      .out(par_reset16_out),
      .done(par_reset16_done)
  );
  
  std_reg #(1) par_done_reg274 (
      .in(par_done_reg274_in),
      .write_en(par_done_reg274_write_en),
      .clk(clk),
      .out(par_done_reg274_out),
      .done(par_done_reg274_done)
  );
  
  std_reg #(1) par_done_reg275 (
      .in(par_done_reg275_in),
      .write_en(par_done_reg275_write_en),
      .clk(clk),
      .out(par_done_reg275_out),
      .done(par_done_reg275_done)
  );
  
  std_reg #(1) par_done_reg276 (
      .in(par_done_reg276_in),
      .write_en(par_done_reg276_write_en),
      .clk(clk),
      .out(par_done_reg276_out),
      .done(par_done_reg276_done)
  );
  
  std_reg #(1) par_done_reg277 (
      .in(par_done_reg277_in),
      .write_en(par_done_reg277_write_en),
      .clk(clk),
      .out(par_done_reg277_out),
      .done(par_done_reg277_done)
  );
  
  std_reg #(1) par_done_reg278 (
      .in(par_done_reg278_in),
      .write_en(par_done_reg278_write_en),
      .clk(clk),
      .out(par_done_reg278_out),
      .done(par_done_reg278_done)
  );
  
  std_reg #(1) par_done_reg279 (
      .in(par_done_reg279_in),
      .write_en(par_done_reg279_write_en),
      .clk(clk),
      .out(par_done_reg279_out),
      .done(par_done_reg279_done)
  );
  
  std_reg #(1) par_done_reg280 (
      .in(par_done_reg280_in),
      .write_en(par_done_reg280_write_en),
      .clk(clk),
      .out(par_done_reg280_out),
      .done(par_done_reg280_done)
  );
  
  std_reg #(1) par_done_reg281 (
      .in(par_done_reg281_in),
      .write_en(par_done_reg281_write_en),
      .clk(clk),
      .out(par_done_reg281_out),
      .done(par_done_reg281_done)
  );
  
  std_reg #(1) par_done_reg282 (
      .in(par_done_reg282_in),
      .write_en(par_done_reg282_write_en),
      .clk(clk),
      .out(par_done_reg282_out),
      .done(par_done_reg282_done)
  );
  
  std_reg #(1) par_done_reg283 (
      .in(par_done_reg283_in),
      .write_en(par_done_reg283_write_en),
      .clk(clk),
      .out(par_done_reg283_out),
      .done(par_done_reg283_done)
  );
  
  std_reg #(1) par_done_reg284 (
      .in(par_done_reg284_in),
      .write_en(par_done_reg284_write_en),
      .clk(clk),
      .out(par_done_reg284_out),
      .done(par_done_reg284_done)
  );
  
  std_reg #(1) par_done_reg285 (
      .in(par_done_reg285_in),
      .write_en(par_done_reg285_write_en),
      .clk(clk),
      .out(par_done_reg285_out),
      .done(par_done_reg285_done)
  );
  
  std_reg #(1) par_done_reg286 (
      .in(par_done_reg286_in),
      .write_en(par_done_reg286_write_en),
      .clk(clk),
      .out(par_done_reg286_out),
      .done(par_done_reg286_done)
  );
  
  std_reg #(1) par_done_reg287 (
      .in(par_done_reg287_in),
      .write_en(par_done_reg287_write_en),
      .clk(clk),
      .out(par_done_reg287_out),
      .done(par_done_reg287_done)
  );
  
  std_reg #(1) par_done_reg288 (
      .in(par_done_reg288_in),
      .write_en(par_done_reg288_write_en),
      .clk(clk),
      .out(par_done_reg288_out),
      .done(par_done_reg288_done)
  );
  
  std_reg #(1) par_done_reg289 (
      .in(par_done_reg289_in),
      .write_en(par_done_reg289_write_en),
      .clk(clk),
      .out(par_done_reg289_out),
      .done(par_done_reg289_done)
  );
  
  std_reg #(1) par_done_reg290 (
      .in(par_done_reg290_in),
      .write_en(par_done_reg290_write_en),
      .clk(clk),
      .out(par_done_reg290_out),
      .done(par_done_reg290_done)
  );
  
  std_reg #(1) par_done_reg291 (
      .in(par_done_reg291_in),
      .write_en(par_done_reg291_write_en),
      .clk(clk),
      .out(par_done_reg291_out),
      .done(par_done_reg291_done)
  );
  
  std_reg #(1) par_done_reg292 (
      .in(par_done_reg292_in),
      .write_en(par_done_reg292_write_en),
      .clk(clk),
      .out(par_done_reg292_out),
      .done(par_done_reg292_done)
  );
  
  std_reg #(1) par_done_reg293 (
      .in(par_done_reg293_in),
      .write_en(par_done_reg293_write_en),
      .clk(clk),
      .out(par_done_reg293_out),
      .done(par_done_reg293_done)
  );
  
  std_reg #(1) par_done_reg294 (
      .in(par_done_reg294_in),
      .write_en(par_done_reg294_write_en),
      .clk(clk),
      .out(par_done_reg294_out),
      .done(par_done_reg294_done)
  );
  
  std_reg #(1) par_done_reg295 (
      .in(par_done_reg295_in),
      .write_en(par_done_reg295_write_en),
      .clk(clk),
      .out(par_done_reg295_out),
      .done(par_done_reg295_done)
  );
  
  std_reg #(1) par_done_reg296 (
      .in(par_done_reg296_in),
      .write_en(par_done_reg296_write_en),
      .clk(clk),
      .out(par_done_reg296_out),
      .done(par_done_reg296_done)
  );
  
  std_reg #(1) par_done_reg297 (
      .in(par_done_reg297_in),
      .write_en(par_done_reg297_write_en),
      .clk(clk),
      .out(par_done_reg297_out),
      .done(par_done_reg297_done)
  );
  
  std_reg #(1) par_done_reg298 (
      .in(par_done_reg298_in),
      .write_en(par_done_reg298_write_en),
      .clk(clk),
      .out(par_done_reg298_out),
      .done(par_done_reg298_done)
  );
  
  std_reg #(1) par_done_reg299 (
      .in(par_done_reg299_in),
      .write_en(par_done_reg299_write_en),
      .clk(clk),
      .out(par_done_reg299_out),
      .done(par_done_reg299_done)
  );
  
  std_reg #(1) par_done_reg300 (
      .in(par_done_reg300_in),
      .write_en(par_done_reg300_write_en),
      .clk(clk),
      .out(par_done_reg300_out),
      .done(par_done_reg300_done)
  );
  
  std_reg #(1) par_done_reg301 (
      .in(par_done_reg301_in),
      .write_en(par_done_reg301_write_en),
      .clk(clk),
      .out(par_done_reg301_out),
      .done(par_done_reg301_done)
  );
  
  std_reg #(1) par_done_reg302 (
      .in(par_done_reg302_in),
      .write_en(par_done_reg302_write_en),
      .clk(clk),
      .out(par_done_reg302_out),
      .done(par_done_reg302_done)
  );
  
  std_reg #(1) par_done_reg303 (
      .in(par_done_reg303_in),
      .write_en(par_done_reg303_write_en),
      .clk(clk),
      .out(par_done_reg303_out),
      .done(par_done_reg303_done)
  );
  
  std_reg #(1) par_done_reg304 (
      .in(par_done_reg304_in),
      .write_en(par_done_reg304_write_en),
      .clk(clk),
      .out(par_done_reg304_out),
      .done(par_done_reg304_done)
  );
  
  std_reg #(1) par_done_reg305 (
      .in(par_done_reg305_in),
      .write_en(par_done_reg305_write_en),
      .clk(clk),
      .out(par_done_reg305_out),
      .done(par_done_reg305_done)
  );
  
  std_reg #(1) par_done_reg306 (
      .in(par_done_reg306_in),
      .write_en(par_done_reg306_write_en),
      .clk(clk),
      .out(par_done_reg306_out),
      .done(par_done_reg306_done)
  );
  
  std_reg #(1) par_done_reg307 (
      .in(par_done_reg307_in),
      .write_en(par_done_reg307_write_en),
      .clk(clk),
      .out(par_done_reg307_out),
      .done(par_done_reg307_done)
  );
  
  std_reg #(1) par_done_reg308 (
      .in(par_done_reg308_in),
      .write_en(par_done_reg308_write_en),
      .clk(clk),
      .out(par_done_reg308_out),
      .done(par_done_reg308_done)
  );
  
  std_reg #(1) par_done_reg309 (
      .in(par_done_reg309_in),
      .write_en(par_done_reg309_write_en),
      .clk(clk),
      .out(par_done_reg309_out),
      .done(par_done_reg309_done)
  );
  
  std_reg #(1) par_reset17 (
      .in(par_reset17_in),
      .write_en(par_reset17_write_en),
      .clk(clk),
      .out(par_reset17_out),
      .done(par_reset17_done)
  );
  
  std_reg #(1) par_done_reg310 (
      .in(par_done_reg310_in),
      .write_en(par_done_reg310_write_en),
      .clk(clk),
      .out(par_done_reg310_out),
      .done(par_done_reg310_done)
  );
  
  std_reg #(1) par_done_reg311 (
      .in(par_done_reg311_in),
      .write_en(par_done_reg311_write_en),
      .clk(clk),
      .out(par_done_reg311_out),
      .done(par_done_reg311_done)
  );
  
  std_reg #(1) par_done_reg312 (
      .in(par_done_reg312_in),
      .write_en(par_done_reg312_write_en),
      .clk(clk),
      .out(par_done_reg312_out),
      .done(par_done_reg312_done)
  );
  
  std_reg #(1) par_done_reg313 (
      .in(par_done_reg313_in),
      .write_en(par_done_reg313_write_en),
      .clk(clk),
      .out(par_done_reg313_out),
      .done(par_done_reg313_done)
  );
  
  std_reg #(1) par_done_reg314 (
      .in(par_done_reg314_in),
      .write_en(par_done_reg314_write_en),
      .clk(clk),
      .out(par_done_reg314_out),
      .done(par_done_reg314_done)
  );
  
  std_reg #(1) par_done_reg315 (
      .in(par_done_reg315_in),
      .write_en(par_done_reg315_write_en),
      .clk(clk),
      .out(par_done_reg315_out),
      .done(par_done_reg315_done)
  );
  
  std_reg #(1) par_done_reg316 (
      .in(par_done_reg316_in),
      .write_en(par_done_reg316_write_en),
      .clk(clk),
      .out(par_done_reg316_out),
      .done(par_done_reg316_done)
  );
  
  std_reg #(1) par_done_reg317 (
      .in(par_done_reg317_in),
      .write_en(par_done_reg317_write_en),
      .clk(clk),
      .out(par_done_reg317_out),
      .done(par_done_reg317_done)
  );
  
  std_reg #(1) par_done_reg318 (
      .in(par_done_reg318_in),
      .write_en(par_done_reg318_write_en),
      .clk(clk),
      .out(par_done_reg318_out),
      .done(par_done_reg318_done)
  );
  
  std_reg #(1) par_done_reg319 (
      .in(par_done_reg319_in),
      .write_en(par_done_reg319_write_en),
      .clk(clk),
      .out(par_done_reg319_out),
      .done(par_done_reg319_done)
  );
  
  std_reg #(1) par_done_reg320 (
      .in(par_done_reg320_in),
      .write_en(par_done_reg320_write_en),
      .clk(clk),
      .out(par_done_reg320_out),
      .done(par_done_reg320_done)
  );
  
  std_reg #(1) par_done_reg321 (
      .in(par_done_reg321_in),
      .write_en(par_done_reg321_write_en),
      .clk(clk),
      .out(par_done_reg321_out),
      .done(par_done_reg321_done)
  );
  
  std_reg #(1) par_done_reg322 (
      .in(par_done_reg322_in),
      .write_en(par_done_reg322_write_en),
      .clk(clk),
      .out(par_done_reg322_out),
      .done(par_done_reg322_done)
  );
  
  std_reg #(1) par_done_reg323 (
      .in(par_done_reg323_in),
      .write_en(par_done_reg323_write_en),
      .clk(clk),
      .out(par_done_reg323_out),
      .done(par_done_reg323_done)
  );
  
  std_reg #(1) par_done_reg324 (
      .in(par_done_reg324_in),
      .write_en(par_done_reg324_write_en),
      .clk(clk),
      .out(par_done_reg324_out),
      .done(par_done_reg324_done)
  );
  
  std_reg #(1) par_done_reg325 (
      .in(par_done_reg325_in),
      .write_en(par_done_reg325_write_en),
      .clk(clk),
      .out(par_done_reg325_out),
      .done(par_done_reg325_done)
  );
  
  std_reg #(1) par_done_reg326 (
      .in(par_done_reg326_in),
      .write_en(par_done_reg326_write_en),
      .clk(clk),
      .out(par_done_reg326_out),
      .done(par_done_reg326_done)
  );
  
  std_reg #(1) par_done_reg327 (
      .in(par_done_reg327_in),
      .write_en(par_done_reg327_write_en),
      .clk(clk),
      .out(par_done_reg327_out),
      .done(par_done_reg327_done)
  );
  
  std_reg #(1) par_done_reg328 (
      .in(par_done_reg328_in),
      .write_en(par_done_reg328_write_en),
      .clk(clk),
      .out(par_done_reg328_out),
      .done(par_done_reg328_done)
  );
  
  std_reg #(1) par_done_reg329 (
      .in(par_done_reg329_in),
      .write_en(par_done_reg329_write_en),
      .clk(clk),
      .out(par_done_reg329_out),
      .done(par_done_reg329_done)
  );
  
  std_reg #(1) par_reset18 (
      .in(par_reset18_in),
      .write_en(par_reset18_write_en),
      .clk(clk),
      .out(par_reset18_out),
      .done(par_reset18_done)
  );
  
  std_reg #(1) par_done_reg330 (
      .in(par_done_reg330_in),
      .write_en(par_done_reg330_write_en),
      .clk(clk),
      .out(par_done_reg330_out),
      .done(par_done_reg330_done)
  );
  
  std_reg #(1) par_done_reg331 (
      .in(par_done_reg331_in),
      .write_en(par_done_reg331_write_en),
      .clk(clk),
      .out(par_done_reg331_out),
      .done(par_done_reg331_done)
  );
  
  std_reg #(1) par_done_reg332 (
      .in(par_done_reg332_in),
      .write_en(par_done_reg332_write_en),
      .clk(clk),
      .out(par_done_reg332_out),
      .done(par_done_reg332_done)
  );
  
  std_reg #(1) par_done_reg333 (
      .in(par_done_reg333_in),
      .write_en(par_done_reg333_write_en),
      .clk(clk),
      .out(par_done_reg333_out),
      .done(par_done_reg333_done)
  );
  
  std_reg #(1) par_done_reg334 (
      .in(par_done_reg334_in),
      .write_en(par_done_reg334_write_en),
      .clk(clk),
      .out(par_done_reg334_out),
      .done(par_done_reg334_done)
  );
  
  std_reg #(1) par_done_reg335 (
      .in(par_done_reg335_in),
      .write_en(par_done_reg335_write_en),
      .clk(clk),
      .out(par_done_reg335_out),
      .done(par_done_reg335_done)
  );
  
  std_reg #(1) par_done_reg336 (
      .in(par_done_reg336_in),
      .write_en(par_done_reg336_write_en),
      .clk(clk),
      .out(par_done_reg336_out),
      .done(par_done_reg336_done)
  );
  
  std_reg #(1) par_done_reg337 (
      .in(par_done_reg337_in),
      .write_en(par_done_reg337_write_en),
      .clk(clk),
      .out(par_done_reg337_out),
      .done(par_done_reg337_done)
  );
  
  std_reg #(1) par_done_reg338 (
      .in(par_done_reg338_in),
      .write_en(par_done_reg338_write_en),
      .clk(clk),
      .out(par_done_reg338_out),
      .done(par_done_reg338_done)
  );
  
  std_reg #(1) par_done_reg339 (
      .in(par_done_reg339_in),
      .write_en(par_done_reg339_write_en),
      .clk(clk),
      .out(par_done_reg339_out),
      .done(par_done_reg339_done)
  );
  
  std_reg #(1) par_done_reg340 (
      .in(par_done_reg340_in),
      .write_en(par_done_reg340_write_en),
      .clk(clk),
      .out(par_done_reg340_out),
      .done(par_done_reg340_done)
  );
  
  std_reg #(1) par_done_reg341 (
      .in(par_done_reg341_in),
      .write_en(par_done_reg341_write_en),
      .clk(clk),
      .out(par_done_reg341_out),
      .done(par_done_reg341_done)
  );
  
  std_reg #(1) par_done_reg342 (
      .in(par_done_reg342_in),
      .write_en(par_done_reg342_write_en),
      .clk(clk),
      .out(par_done_reg342_out),
      .done(par_done_reg342_done)
  );
  
  std_reg #(1) par_done_reg343 (
      .in(par_done_reg343_in),
      .write_en(par_done_reg343_write_en),
      .clk(clk),
      .out(par_done_reg343_out),
      .done(par_done_reg343_done)
  );
  
  std_reg #(1) par_done_reg344 (
      .in(par_done_reg344_in),
      .write_en(par_done_reg344_write_en),
      .clk(clk),
      .out(par_done_reg344_out),
      .done(par_done_reg344_done)
  );
  
  std_reg #(1) par_done_reg345 (
      .in(par_done_reg345_in),
      .write_en(par_done_reg345_write_en),
      .clk(clk),
      .out(par_done_reg345_out),
      .done(par_done_reg345_done)
  );
  
  std_reg #(1) par_done_reg346 (
      .in(par_done_reg346_in),
      .write_en(par_done_reg346_write_en),
      .clk(clk),
      .out(par_done_reg346_out),
      .done(par_done_reg346_done)
  );
  
  std_reg #(1) par_done_reg347 (
      .in(par_done_reg347_in),
      .write_en(par_done_reg347_write_en),
      .clk(clk),
      .out(par_done_reg347_out),
      .done(par_done_reg347_done)
  );
  
  std_reg #(1) par_done_reg348 (
      .in(par_done_reg348_in),
      .write_en(par_done_reg348_write_en),
      .clk(clk),
      .out(par_done_reg348_out),
      .done(par_done_reg348_done)
  );
  
  std_reg #(1) par_done_reg349 (
      .in(par_done_reg349_in),
      .write_en(par_done_reg349_write_en),
      .clk(clk),
      .out(par_done_reg349_out),
      .done(par_done_reg349_done)
  );
  
  std_reg #(1) par_done_reg350 (
      .in(par_done_reg350_in),
      .write_en(par_done_reg350_write_en),
      .clk(clk),
      .out(par_done_reg350_out),
      .done(par_done_reg350_done)
  );
  
  std_reg #(1) par_done_reg351 (
      .in(par_done_reg351_in),
      .write_en(par_done_reg351_write_en),
      .clk(clk),
      .out(par_done_reg351_out),
      .done(par_done_reg351_done)
  );
  
  std_reg #(1) par_done_reg352 (
      .in(par_done_reg352_in),
      .write_en(par_done_reg352_write_en),
      .clk(clk),
      .out(par_done_reg352_out),
      .done(par_done_reg352_done)
  );
  
  std_reg #(1) par_done_reg353 (
      .in(par_done_reg353_in),
      .write_en(par_done_reg353_write_en),
      .clk(clk),
      .out(par_done_reg353_out),
      .done(par_done_reg353_done)
  );
  
  std_reg #(1) par_done_reg354 (
      .in(par_done_reg354_in),
      .write_en(par_done_reg354_write_en),
      .clk(clk),
      .out(par_done_reg354_out),
      .done(par_done_reg354_done)
  );
  
  std_reg #(1) par_done_reg355 (
      .in(par_done_reg355_in),
      .write_en(par_done_reg355_write_en),
      .clk(clk),
      .out(par_done_reg355_out),
      .done(par_done_reg355_done)
  );
  
  std_reg #(1) par_done_reg356 (
      .in(par_done_reg356_in),
      .write_en(par_done_reg356_write_en),
      .clk(clk),
      .out(par_done_reg356_out),
      .done(par_done_reg356_done)
  );
  
  std_reg #(1) par_done_reg357 (
      .in(par_done_reg357_in),
      .write_en(par_done_reg357_write_en),
      .clk(clk),
      .out(par_done_reg357_out),
      .done(par_done_reg357_done)
  );
  
  std_reg #(1) par_done_reg358 (
      .in(par_done_reg358_in),
      .write_en(par_done_reg358_write_en),
      .clk(clk),
      .out(par_done_reg358_out),
      .done(par_done_reg358_done)
  );
  
  std_reg #(1) par_done_reg359 (
      .in(par_done_reg359_in),
      .write_en(par_done_reg359_write_en),
      .clk(clk),
      .out(par_done_reg359_out),
      .done(par_done_reg359_done)
  );
  
  std_reg #(1) par_reset19 (
      .in(par_reset19_in),
      .write_en(par_reset19_write_en),
      .clk(clk),
      .out(par_reset19_out),
      .done(par_reset19_done)
  );
  
  std_reg #(1) par_done_reg360 (
      .in(par_done_reg360_in),
      .write_en(par_done_reg360_write_en),
      .clk(clk),
      .out(par_done_reg360_out),
      .done(par_done_reg360_done)
  );
  
  std_reg #(1) par_done_reg361 (
      .in(par_done_reg361_in),
      .write_en(par_done_reg361_write_en),
      .clk(clk),
      .out(par_done_reg361_out),
      .done(par_done_reg361_done)
  );
  
  std_reg #(1) par_done_reg362 (
      .in(par_done_reg362_in),
      .write_en(par_done_reg362_write_en),
      .clk(clk),
      .out(par_done_reg362_out),
      .done(par_done_reg362_done)
  );
  
  std_reg #(1) par_done_reg363 (
      .in(par_done_reg363_in),
      .write_en(par_done_reg363_write_en),
      .clk(clk),
      .out(par_done_reg363_out),
      .done(par_done_reg363_done)
  );
  
  std_reg #(1) par_done_reg364 (
      .in(par_done_reg364_in),
      .write_en(par_done_reg364_write_en),
      .clk(clk),
      .out(par_done_reg364_out),
      .done(par_done_reg364_done)
  );
  
  std_reg #(1) par_done_reg365 (
      .in(par_done_reg365_in),
      .write_en(par_done_reg365_write_en),
      .clk(clk),
      .out(par_done_reg365_out),
      .done(par_done_reg365_done)
  );
  
  std_reg #(1) par_done_reg366 (
      .in(par_done_reg366_in),
      .write_en(par_done_reg366_write_en),
      .clk(clk),
      .out(par_done_reg366_out),
      .done(par_done_reg366_done)
  );
  
  std_reg #(1) par_done_reg367 (
      .in(par_done_reg367_in),
      .write_en(par_done_reg367_write_en),
      .clk(clk),
      .out(par_done_reg367_out),
      .done(par_done_reg367_done)
  );
  
  std_reg #(1) par_done_reg368 (
      .in(par_done_reg368_in),
      .write_en(par_done_reg368_write_en),
      .clk(clk),
      .out(par_done_reg368_out),
      .done(par_done_reg368_done)
  );
  
  std_reg #(1) par_done_reg369 (
      .in(par_done_reg369_in),
      .write_en(par_done_reg369_write_en),
      .clk(clk),
      .out(par_done_reg369_out),
      .done(par_done_reg369_done)
  );
  
  std_reg #(1) par_done_reg370 (
      .in(par_done_reg370_in),
      .write_en(par_done_reg370_write_en),
      .clk(clk),
      .out(par_done_reg370_out),
      .done(par_done_reg370_done)
  );
  
  std_reg #(1) par_done_reg371 (
      .in(par_done_reg371_in),
      .write_en(par_done_reg371_write_en),
      .clk(clk),
      .out(par_done_reg371_out),
      .done(par_done_reg371_done)
  );
  
  std_reg #(1) par_done_reg372 (
      .in(par_done_reg372_in),
      .write_en(par_done_reg372_write_en),
      .clk(clk),
      .out(par_done_reg372_out),
      .done(par_done_reg372_done)
  );
  
  std_reg #(1) par_done_reg373 (
      .in(par_done_reg373_in),
      .write_en(par_done_reg373_write_en),
      .clk(clk),
      .out(par_done_reg373_out),
      .done(par_done_reg373_done)
  );
  
  std_reg #(1) par_done_reg374 (
      .in(par_done_reg374_in),
      .write_en(par_done_reg374_write_en),
      .clk(clk),
      .out(par_done_reg374_out),
      .done(par_done_reg374_done)
  );
  
  std_reg #(1) par_reset20 (
      .in(par_reset20_in),
      .write_en(par_reset20_write_en),
      .clk(clk),
      .out(par_reset20_out),
      .done(par_reset20_done)
  );
  
  std_reg #(1) par_done_reg375 (
      .in(par_done_reg375_in),
      .write_en(par_done_reg375_write_en),
      .clk(clk),
      .out(par_done_reg375_out),
      .done(par_done_reg375_done)
  );
  
  std_reg #(1) par_done_reg376 (
      .in(par_done_reg376_in),
      .write_en(par_done_reg376_write_en),
      .clk(clk),
      .out(par_done_reg376_out),
      .done(par_done_reg376_done)
  );
  
  std_reg #(1) par_done_reg377 (
      .in(par_done_reg377_in),
      .write_en(par_done_reg377_write_en),
      .clk(clk),
      .out(par_done_reg377_out),
      .done(par_done_reg377_done)
  );
  
  std_reg #(1) par_done_reg378 (
      .in(par_done_reg378_in),
      .write_en(par_done_reg378_write_en),
      .clk(clk),
      .out(par_done_reg378_out),
      .done(par_done_reg378_done)
  );
  
  std_reg #(1) par_done_reg379 (
      .in(par_done_reg379_in),
      .write_en(par_done_reg379_write_en),
      .clk(clk),
      .out(par_done_reg379_out),
      .done(par_done_reg379_done)
  );
  
  std_reg #(1) par_done_reg380 (
      .in(par_done_reg380_in),
      .write_en(par_done_reg380_write_en),
      .clk(clk),
      .out(par_done_reg380_out),
      .done(par_done_reg380_done)
  );
  
  std_reg #(1) par_done_reg381 (
      .in(par_done_reg381_in),
      .write_en(par_done_reg381_write_en),
      .clk(clk),
      .out(par_done_reg381_out),
      .done(par_done_reg381_done)
  );
  
  std_reg #(1) par_done_reg382 (
      .in(par_done_reg382_in),
      .write_en(par_done_reg382_write_en),
      .clk(clk),
      .out(par_done_reg382_out),
      .done(par_done_reg382_done)
  );
  
  std_reg #(1) par_done_reg383 (
      .in(par_done_reg383_in),
      .write_en(par_done_reg383_write_en),
      .clk(clk),
      .out(par_done_reg383_out),
      .done(par_done_reg383_done)
  );
  
  std_reg #(1) par_done_reg384 (
      .in(par_done_reg384_in),
      .write_en(par_done_reg384_write_en),
      .clk(clk),
      .out(par_done_reg384_out),
      .done(par_done_reg384_done)
  );
  
  std_reg #(1) par_done_reg385 (
      .in(par_done_reg385_in),
      .write_en(par_done_reg385_write_en),
      .clk(clk),
      .out(par_done_reg385_out),
      .done(par_done_reg385_done)
  );
  
  std_reg #(1) par_done_reg386 (
      .in(par_done_reg386_in),
      .write_en(par_done_reg386_write_en),
      .clk(clk),
      .out(par_done_reg386_out),
      .done(par_done_reg386_done)
  );
  
  std_reg #(1) par_done_reg387 (
      .in(par_done_reg387_in),
      .write_en(par_done_reg387_write_en),
      .clk(clk),
      .out(par_done_reg387_out),
      .done(par_done_reg387_done)
  );
  
  std_reg #(1) par_done_reg388 (
      .in(par_done_reg388_in),
      .write_en(par_done_reg388_write_en),
      .clk(clk),
      .out(par_done_reg388_out),
      .done(par_done_reg388_done)
  );
  
  std_reg #(1) par_done_reg389 (
      .in(par_done_reg389_in),
      .write_en(par_done_reg389_write_en),
      .clk(clk),
      .out(par_done_reg389_out),
      .done(par_done_reg389_done)
  );
  
  std_reg #(1) par_done_reg390 (
      .in(par_done_reg390_in),
      .write_en(par_done_reg390_write_en),
      .clk(clk),
      .out(par_done_reg390_out),
      .done(par_done_reg390_done)
  );
  
  std_reg #(1) par_done_reg391 (
      .in(par_done_reg391_in),
      .write_en(par_done_reg391_write_en),
      .clk(clk),
      .out(par_done_reg391_out),
      .done(par_done_reg391_done)
  );
  
  std_reg #(1) par_done_reg392 (
      .in(par_done_reg392_in),
      .write_en(par_done_reg392_write_en),
      .clk(clk),
      .out(par_done_reg392_out),
      .done(par_done_reg392_done)
  );
  
  std_reg #(1) par_done_reg393 (
      .in(par_done_reg393_in),
      .write_en(par_done_reg393_write_en),
      .clk(clk),
      .out(par_done_reg393_out),
      .done(par_done_reg393_done)
  );
  
  std_reg #(1) par_done_reg394 (
      .in(par_done_reg394_in),
      .write_en(par_done_reg394_write_en),
      .clk(clk),
      .out(par_done_reg394_out),
      .done(par_done_reg394_done)
  );
  
  std_reg #(1) par_reset21 (
      .in(par_reset21_in),
      .write_en(par_reset21_write_en),
      .clk(clk),
      .out(par_reset21_out),
      .done(par_reset21_done)
  );
  
  std_reg #(1) par_done_reg395 (
      .in(par_done_reg395_in),
      .write_en(par_done_reg395_write_en),
      .clk(clk),
      .out(par_done_reg395_out),
      .done(par_done_reg395_done)
  );
  
  std_reg #(1) par_done_reg396 (
      .in(par_done_reg396_in),
      .write_en(par_done_reg396_write_en),
      .clk(clk),
      .out(par_done_reg396_out),
      .done(par_done_reg396_done)
  );
  
  std_reg #(1) par_done_reg397 (
      .in(par_done_reg397_in),
      .write_en(par_done_reg397_write_en),
      .clk(clk),
      .out(par_done_reg397_out),
      .done(par_done_reg397_done)
  );
  
  std_reg #(1) par_done_reg398 (
      .in(par_done_reg398_in),
      .write_en(par_done_reg398_write_en),
      .clk(clk),
      .out(par_done_reg398_out),
      .done(par_done_reg398_done)
  );
  
  std_reg #(1) par_done_reg399 (
      .in(par_done_reg399_in),
      .write_en(par_done_reg399_write_en),
      .clk(clk),
      .out(par_done_reg399_out),
      .done(par_done_reg399_done)
  );
  
  std_reg #(1) par_done_reg400 (
      .in(par_done_reg400_in),
      .write_en(par_done_reg400_write_en),
      .clk(clk),
      .out(par_done_reg400_out),
      .done(par_done_reg400_done)
  );
  
  std_reg #(1) par_done_reg401 (
      .in(par_done_reg401_in),
      .write_en(par_done_reg401_write_en),
      .clk(clk),
      .out(par_done_reg401_out),
      .done(par_done_reg401_done)
  );
  
  std_reg #(1) par_done_reg402 (
      .in(par_done_reg402_in),
      .write_en(par_done_reg402_write_en),
      .clk(clk),
      .out(par_done_reg402_out),
      .done(par_done_reg402_done)
  );
  
  std_reg #(1) par_done_reg403 (
      .in(par_done_reg403_in),
      .write_en(par_done_reg403_write_en),
      .clk(clk),
      .out(par_done_reg403_out),
      .done(par_done_reg403_done)
  );
  
  std_reg #(1) par_done_reg404 (
      .in(par_done_reg404_in),
      .write_en(par_done_reg404_write_en),
      .clk(clk),
      .out(par_done_reg404_out),
      .done(par_done_reg404_done)
  );
  
  std_reg #(1) par_reset22 (
      .in(par_reset22_in),
      .write_en(par_reset22_write_en),
      .clk(clk),
      .out(par_reset22_out),
      .done(par_reset22_done)
  );
  
  std_reg #(1) par_done_reg405 (
      .in(par_done_reg405_in),
      .write_en(par_done_reg405_write_en),
      .clk(clk),
      .out(par_done_reg405_out),
      .done(par_done_reg405_done)
  );
  
  std_reg #(1) par_done_reg406 (
      .in(par_done_reg406_in),
      .write_en(par_done_reg406_write_en),
      .clk(clk),
      .out(par_done_reg406_out),
      .done(par_done_reg406_done)
  );
  
  std_reg #(1) par_done_reg407 (
      .in(par_done_reg407_in),
      .write_en(par_done_reg407_write_en),
      .clk(clk),
      .out(par_done_reg407_out),
      .done(par_done_reg407_done)
  );
  
  std_reg #(1) par_done_reg408 (
      .in(par_done_reg408_in),
      .write_en(par_done_reg408_write_en),
      .clk(clk),
      .out(par_done_reg408_out),
      .done(par_done_reg408_done)
  );
  
  std_reg #(1) par_done_reg409 (
      .in(par_done_reg409_in),
      .write_en(par_done_reg409_write_en),
      .clk(clk),
      .out(par_done_reg409_out),
      .done(par_done_reg409_done)
  );
  
  std_reg #(1) par_done_reg410 (
      .in(par_done_reg410_in),
      .write_en(par_done_reg410_write_en),
      .clk(clk),
      .out(par_done_reg410_out),
      .done(par_done_reg410_done)
  );
  
  std_reg #(1) par_done_reg411 (
      .in(par_done_reg411_in),
      .write_en(par_done_reg411_write_en),
      .clk(clk),
      .out(par_done_reg411_out),
      .done(par_done_reg411_done)
  );
  
  std_reg #(1) par_done_reg412 (
      .in(par_done_reg412_in),
      .write_en(par_done_reg412_write_en),
      .clk(clk),
      .out(par_done_reg412_out),
      .done(par_done_reg412_done)
  );
  
  std_reg #(1) par_done_reg413 (
      .in(par_done_reg413_in),
      .write_en(par_done_reg413_write_en),
      .clk(clk),
      .out(par_done_reg413_out),
      .done(par_done_reg413_done)
  );
  
  std_reg #(1) par_done_reg414 (
      .in(par_done_reg414_in),
      .write_en(par_done_reg414_write_en),
      .clk(clk),
      .out(par_done_reg414_out),
      .done(par_done_reg414_done)
  );
  
  std_reg #(1) par_done_reg415 (
      .in(par_done_reg415_in),
      .write_en(par_done_reg415_write_en),
      .clk(clk),
      .out(par_done_reg415_out),
      .done(par_done_reg415_done)
  );
  
  std_reg #(1) par_done_reg416 (
      .in(par_done_reg416_in),
      .write_en(par_done_reg416_write_en),
      .clk(clk),
      .out(par_done_reg416_out),
      .done(par_done_reg416_done)
  );
  
  std_reg #(1) par_reset23 (
      .in(par_reset23_in),
      .write_en(par_reset23_write_en),
      .clk(clk),
      .out(par_reset23_out),
      .done(par_reset23_done)
  );
  
  std_reg #(1) par_done_reg417 (
      .in(par_done_reg417_in),
      .write_en(par_done_reg417_write_en),
      .clk(clk),
      .out(par_done_reg417_out),
      .done(par_done_reg417_done)
  );
  
  std_reg #(1) par_done_reg418 (
      .in(par_done_reg418_in),
      .write_en(par_done_reg418_write_en),
      .clk(clk),
      .out(par_done_reg418_out),
      .done(par_done_reg418_done)
  );
  
  std_reg #(1) par_done_reg419 (
      .in(par_done_reg419_in),
      .write_en(par_done_reg419_write_en),
      .clk(clk),
      .out(par_done_reg419_out),
      .done(par_done_reg419_done)
  );
  
  std_reg #(1) par_done_reg420 (
      .in(par_done_reg420_in),
      .write_en(par_done_reg420_write_en),
      .clk(clk),
      .out(par_done_reg420_out),
      .done(par_done_reg420_done)
  );
  
  std_reg #(1) par_done_reg421 (
      .in(par_done_reg421_in),
      .write_en(par_done_reg421_write_en),
      .clk(clk),
      .out(par_done_reg421_out),
      .done(par_done_reg421_done)
  );
  
  std_reg #(1) par_done_reg422 (
      .in(par_done_reg422_in),
      .write_en(par_done_reg422_write_en),
      .clk(clk),
      .out(par_done_reg422_out),
      .done(par_done_reg422_done)
  );
  
  std_reg #(1) par_reset24 (
      .in(par_reset24_in),
      .write_en(par_reset24_write_en),
      .clk(clk),
      .out(par_reset24_out),
      .done(par_reset24_done)
  );
  
  std_reg #(1) par_done_reg423 (
      .in(par_done_reg423_in),
      .write_en(par_done_reg423_write_en),
      .clk(clk),
      .out(par_done_reg423_out),
      .done(par_done_reg423_done)
  );
  
  std_reg #(1) par_done_reg424 (
      .in(par_done_reg424_in),
      .write_en(par_done_reg424_write_en),
      .clk(clk),
      .out(par_done_reg424_out),
      .done(par_done_reg424_done)
  );
  
  std_reg #(1) par_done_reg425 (
      .in(par_done_reg425_in),
      .write_en(par_done_reg425_write_en),
      .clk(clk),
      .out(par_done_reg425_out),
      .done(par_done_reg425_done)
  );
  
  std_reg #(1) par_done_reg426 (
      .in(par_done_reg426_in),
      .write_en(par_done_reg426_write_en),
      .clk(clk),
      .out(par_done_reg426_out),
      .done(par_done_reg426_done)
  );
  
  std_reg #(1) par_done_reg427 (
      .in(par_done_reg427_in),
      .write_en(par_done_reg427_write_en),
      .clk(clk),
      .out(par_done_reg427_out),
      .done(par_done_reg427_done)
  );
  
  std_reg #(1) par_done_reg428 (
      .in(par_done_reg428_in),
      .write_en(par_done_reg428_write_en),
      .clk(clk),
      .out(par_done_reg428_out),
      .done(par_done_reg428_done)
  );
  
  std_reg #(1) par_reset25 (
      .in(par_reset25_in),
      .write_en(par_reset25_write_en),
      .clk(clk),
      .out(par_reset25_out),
      .done(par_reset25_done)
  );
  
  std_reg #(1) par_done_reg429 (
      .in(par_done_reg429_in),
      .write_en(par_done_reg429_write_en),
      .clk(clk),
      .out(par_done_reg429_out),
      .done(par_done_reg429_done)
  );
  
  std_reg #(1) par_done_reg430 (
      .in(par_done_reg430_in),
      .write_en(par_done_reg430_write_en),
      .clk(clk),
      .out(par_done_reg430_out),
      .done(par_done_reg430_done)
  );
  
  std_reg #(1) par_done_reg431 (
      .in(par_done_reg431_in),
      .write_en(par_done_reg431_write_en),
      .clk(clk),
      .out(par_done_reg431_out),
      .done(par_done_reg431_done)
  );
  
  std_reg #(1) par_reset26 (
      .in(par_reset26_in),
      .write_en(par_reset26_write_en),
      .clk(clk),
      .out(par_reset26_out),
      .done(par_reset26_done)
  );
  
  std_reg #(1) par_done_reg432 (
      .in(par_done_reg432_in),
      .write_en(par_done_reg432_write_en),
      .clk(clk),
      .out(par_done_reg432_out),
      .done(par_done_reg432_done)
  );
  
  std_reg #(1) par_done_reg433 (
      .in(par_done_reg433_in),
      .write_en(par_done_reg433_write_en),
      .clk(clk),
      .out(par_done_reg433_out),
      .done(par_done_reg433_done)
  );
  
  std_reg #(1) par_reset27 (
      .in(par_reset27_in),
      .write_en(par_reset27_write_en),
      .clk(clk),
      .out(par_reset27_out),
      .done(par_reset27_done)
  );
  
  std_reg #(1) par_done_reg434 (
      .in(par_done_reg434_in),
      .write_en(par_done_reg434_write_en),
      .clk(clk),
      .out(par_done_reg434_out),
      .done(par_done_reg434_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign done = (fsm0_out == 32'd53) ? 1'd1 : '0;
  assign out_mem_addr0 = (fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go) ? 3'd4 : (fsm0_out == 32'd43 & !out_mem_done & go | fsm0_out == 32'd44 & !out_mem_done & go | fsm0_out == 32'd45 & !out_mem_done & go | fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go) ? 3'd3 : (fsm0_out == 32'd38 & !out_mem_done & go | fsm0_out == 32'd39 & !out_mem_done & go | fsm0_out == 32'd40 & !out_mem_done & go | fsm0_out == 32'd41 & !out_mem_done & go | fsm0_out == 32'd42 & !out_mem_done & go) ? 3'd2 : (fsm0_out == 32'd28 & !out_mem_done & go | fsm0_out == 32'd29 & !out_mem_done & go | fsm0_out == 32'd30 & !out_mem_done & go | fsm0_out == 32'd31 & !out_mem_done & go | fsm0_out == 32'd32 & !out_mem_done & go) ? 3'd0 : (fsm0_out == 32'd33 & !out_mem_done & go | fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go) ? 3'd1 : '0;
  assign out_mem_addr1 = (fsm0_out == 32'd32 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go | fsm0_out == 32'd42 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go) ? 3'd4 : (fsm0_out == 32'd31 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd41 & !out_mem_done & go | fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go) ? 3'd3 : (fsm0_out == 32'd30 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd40 & !out_mem_done & go | fsm0_out == 32'd45 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go) ? 3'd2 : (fsm0_out == 32'd28 & !out_mem_done & go | fsm0_out == 32'd33 & !out_mem_done & go | fsm0_out == 32'd38 & !out_mem_done & go | fsm0_out == 32'd43 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go) ? 3'd0 : (fsm0_out == 32'd29 & !out_mem_done & go | fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd39 & !out_mem_done & go | fsm0_out == 32'd44 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go) ? 3'd1 : '0;
  assign out_mem_write_data = (fsm0_out == 32'd52 & !out_mem_done & go) ? pe_44_out : (fsm0_out == 32'd51 & !out_mem_done & go) ? pe_43_out : (fsm0_out == 32'd50 & !out_mem_done & go) ? pe_42_out : (fsm0_out == 32'd49 & !out_mem_done & go) ? pe_41_out : (fsm0_out == 32'd48 & !out_mem_done & go) ? pe_40_out : (fsm0_out == 32'd47 & !out_mem_done & go) ? pe_34_out : (fsm0_out == 32'd46 & !out_mem_done & go) ? pe_33_out : (fsm0_out == 32'd45 & !out_mem_done & go) ? pe_32_out : (fsm0_out == 32'd44 & !out_mem_done & go) ? pe_31_out : (fsm0_out == 32'd43 & !out_mem_done & go) ? pe_30_out : (fsm0_out == 32'd42 & !out_mem_done & go) ? pe_24_out : (fsm0_out == 32'd41 & !out_mem_done & go) ? pe_23_out : (fsm0_out == 32'd40 & !out_mem_done & go) ? pe_22_out : (fsm0_out == 32'd39 & !out_mem_done & go) ? pe_21_out : (fsm0_out == 32'd38 & !out_mem_done & go) ? pe_20_out : (fsm0_out == 32'd37 & !out_mem_done & go) ? pe_14_out : (fsm0_out == 32'd36 & !out_mem_done & go) ? pe_13_out : (fsm0_out == 32'd35 & !out_mem_done & go) ? pe_12_out : (fsm0_out == 32'd34 & !out_mem_done & go) ? pe_11_out : (fsm0_out == 32'd33 & !out_mem_done & go) ? pe_10_out : (fsm0_out == 32'd32 & !out_mem_done & go) ? pe_04_out : (fsm0_out == 32'd31 & !out_mem_done & go) ? pe_03_out : (fsm0_out == 32'd30 & !out_mem_done & go) ? pe_02_out : (fsm0_out == 32'd29 & !out_mem_done & go) ? pe_01_out : (fsm0_out == 32'd28 & !out_mem_done & go) ? pe_00_out : '0;
  assign out_mem_write_en = (fsm0_out == 32'd28 & !out_mem_done & go | fsm0_out == 32'd29 & !out_mem_done & go | fsm0_out == 32'd30 & !out_mem_done & go | fsm0_out == 32'd31 & !out_mem_done & go | fsm0_out == 32'd32 & !out_mem_done & go | fsm0_out == 32'd33 & !out_mem_done & go | fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go | fsm0_out == 32'd38 & !out_mem_done & go | fsm0_out == 32'd39 & !out_mem_done & go | fsm0_out == 32'd40 & !out_mem_done & go | fsm0_out == 32'd41 & !out_mem_done & go | fsm0_out == 32'd42 & !out_mem_done & go | fsm0_out == 32'd43 & !out_mem_done & go | fsm0_out == 32'd44 & !out_mem_done & go | fsm0_out == 32'd45 & !out_mem_done & go | fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go) ? 1'd1 : '0;
  assign left_44_read_in = (!(par_done_reg359_out | left_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg394_out | left_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg416_out | left_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg428_out | left_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg433_out | left_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_43_write_out : '0;
  assign left_44_read_write_en = (!(par_done_reg359_out | left_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg394_out | left_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg416_out | left_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg428_out | left_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg433_out | left_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_44_read_in = (!(par_done_reg344_out | top_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg384_out | top_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg410_out | top_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg425_out | top_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg432_out | top_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_34_write_out : '0;
  assign top_44_read_write_en = (!(par_done_reg344_out | top_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg384_out | top_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg410_out | top_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg425_out | top_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg432_out | top_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_44_top = (!(par_done_reg374_out | pe_44_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg404_out | pe_44_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg422_out | pe_44_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg431_out | pe_44_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg434_out | pe_44_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_44_read_out : '0;
  assign pe_44_left = (!(par_done_reg374_out | pe_44_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg404_out | pe_44_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg422_out | pe_44_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg431_out | pe_44_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg434_out | pe_44_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_44_read_out : '0;
  assign pe_44_go = (!pe_44_done & (!(par_done_reg374_out | pe_44_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg404_out | pe_44_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg422_out | pe_44_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg431_out | pe_44_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg434_out | pe_44_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_43_write_in = (pe_43_done & (!(par_done_reg329_out | right_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg373_out | right_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg403_out | right_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg421_out | right_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg430_out | right_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_43_right : '0;
  assign right_43_write_write_en = (pe_43_done & (!(par_done_reg329_out | right_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg373_out | right_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg403_out | right_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg421_out | right_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg430_out | right_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_43_read_in = (!(par_done_reg309_out | left_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg358_out | left_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg393_out | left_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg415_out | left_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg427_out | left_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_42_write_out : '0;
  assign left_43_read_write_en = (!(par_done_reg309_out | left_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg358_out | left_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg393_out | left_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg415_out | left_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg427_out | left_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_43_read_in = (!(par_done_reg291_out | top_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg343_out | top_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg383_out | top_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg409_out | top_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg424_out | top_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_33_write_out : '0;
  assign top_43_read_write_en = (!(par_done_reg291_out | top_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg343_out | top_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg383_out | top_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg409_out | top_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg424_out | top_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_43_top = (!(par_done_reg329_out | right_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg373_out | right_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg403_out | right_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg421_out | right_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg430_out | right_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_43_read_out : '0;
  assign pe_43_left = (!(par_done_reg329_out | right_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg373_out | right_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg403_out | right_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg421_out | right_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg430_out | right_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_43_read_out : '0;
  assign pe_43_go = (!pe_43_done & (!(par_done_reg329_out | right_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg373_out | right_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg403_out | right_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg421_out | right_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg430_out | right_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_42_write_in = (pe_42_done & (!(par_done_reg273_out | right_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg328_out | right_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg372_out | right_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg402_out | right_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg420_out | right_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_42_right : '0;
  assign right_42_write_write_en = (pe_42_done & (!(par_done_reg273_out | right_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg328_out | right_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg372_out | right_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg402_out | right_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg420_out | right_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_42_read_in = (!(par_done_reg250_out | left_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg308_out | left_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg357_out | left_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg392_out | left_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg414_out | left_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_41_write_out : '0;
  assign left_42_read_write_en = (!(par_done_reg250_out | left_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg308_out | left_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg357_out | left_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg392_out | left_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg414_out | left_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_42_read_in = (!(par_done_reg231_out | top_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg290_out | top_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg342_out | top_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg382_out | top_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg408_out | top_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_32_write_out : '0;
  assign top_42_read_write_en = (!(par_done_reg231_out | top_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg290_out | top_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg342_out | top_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg382_out | top_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg408_out | top_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_42_top = (!(par_done_reg273_out | right_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg328_out | right_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg372_out | right_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg402_out | right_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg420_out | right_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_42_read_out : '0;
  assign pe_42_left = (!(par_done_reg273_out | right_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg328_out | right_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg372_out | right_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg402_out | right_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg420_out | right_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_42_read_out : '0;
  assign pe_42_go = (!pe_42_done & (!(par_done_reg273_out | right_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg328_out | right_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg372_out | right_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg402_out | right_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg420_out | right_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_41_write_in = (pe_41_done & (!(par_done_reg212_out | right_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg272_out | right_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg327_out | right_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg371_out | right_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg401_out | right_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_41_right : '0;
  assign right_41_write_write_en = (pe_41_done & (!(par_done_reg212_out | right_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg272_out | right_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg327_out | right_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg371_out | right_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg401_out | right_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_41_read_in = (!(par_done_reg188_out | left_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg249_out | left_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg307_out | left_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg356_out | left_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg391_out | left_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_40_write_out : '0;
  assign left_41_read_write_en = (!(par_done_reg188_out | left_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg249_out | left_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg307_out | left_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg356_out | left_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg391_out | left_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_41_read_in = (!(par_done_reg170_out | top_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg230_out | top_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg289_out | top_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg341_out | top_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg381_out | top_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_31_write_out : '0;
  assign top_41_read_write_en = (!(par_done_reg170_out | top_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg230_out | top_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg289_out | top_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg341_out | top_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg381_out | top_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_41_top = (!(par_done_reg212_out | right_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg272_out | right_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg327_out | right_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg371_out | right_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg401_out | right_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_41_read_out : '0;
  assign pe_41_left = (!(par_done_reg212_out | right_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg272_out | right_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg327_out | right_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg371_out | right_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg401_out | right_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_41_read_out : '0;
  assign pe_41_go = (!pe_41_done & (!(par_done_reg212_out | right_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg272_out | right_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg327_out | right_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg371_out | right_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg401_out | right_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_40_write_in = (pe_40_done & (!(par_done_reg152_out | right_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg271_out | right_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg326_out | right_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg370_out | right_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_40_right : '0;
  assign right_40_write_write_en = (pe_40_done & (!(par_done_reg152_out | right_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg271_out | right_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg326_out | right_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg370_out | right_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_40_read_in = (!(par_done_reg129_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg306_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg355_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? l4_read_data : '0;
  assign left_40_read_write_en = (!(par_done_reg129_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg306_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg355_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_40_read_in = (!(par_done_reg114_out | top_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg169_out | top_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg229_out | top_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg288_out | top_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg340_out | top_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_30_write_out : '0;
  assign top_40_read_write_en = (!(par_done_reg114_out | top_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg169_out | top_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg229_out | top_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg288_out | top_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg340_out | top_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_40_top = (!(par_done_reg152_out | right_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg271_out | right_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg326_out | right_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg370_out | right_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_40_read_out : '0;
  assign pe_40_left = (!(par_done_reg152_out | right_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg271_out | right_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg326_out | right_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg370_out | right_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_40_read_out : '0;
  assign pe_40_go = (!pe_40_done & (!(par_done_reg152_out | right_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg271_out | right_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg326_out | right_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg370_out | right_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_34_write_in = (pe_34_done & (!(par_done_reg325_out | down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg369_out | down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg400_out | down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg419_out | down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg429_out | down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_34_down : '0;
  assign down_34_write_write_en = (pe_34_done & (!(par_done_reg325_out | down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg369_out | down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg400_out | down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg419_out | down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg429_out | down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_34_read_in = (!(par_done_reg305_out | left_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg354_out | left_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg390_out | left_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg413_out | left_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg426_out | left_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_33_write_out : '0;
  assign left_34_read_write_en = (!(par_done_reg305_out | left_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg354_out | left_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg390_out | left_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg413_out | left_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg426_out | left_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_34_read_in = (!(par_done_reg287_out | top_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg339_out | top_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg380_out | top_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg407_out | top_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg423_out | top_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_24_write_out : '0;
  assign top_34_read_write_en = (!(par_done_reg287_out | top_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg339_out | top_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg380_out | top_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg407_out | top_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg423_out | top_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_34_top = (!(par_done_reg325_out | down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg369_out | down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg400_out | down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg419_out | down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg429_out | down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_34_read_out : '0;
  assign pe_34_left = (!(par_done_reg325_out | down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg369_out | down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg400_out | down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg419_out | down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg429_out | down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_34_read_out : '0;
  assign pe_34_go = (!pe_34_done & (!(par_done_reg325_out | down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg369_out | down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg400_out | down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg419_out | down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg429_out | down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_33_write_in = (pe_33_done & (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_33_down : '0;
  assign down_33_write_write_en = (pe_33_done & (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_33_write_in = (pe_33_done & (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_33_right : '0;
  assign right_33_write_write_en = (pe_33_done & (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_33_read_in = (!(par_done_reg247_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg304_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg353_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg389_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg412_out | left_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_32_write_out : '0;
  assign left_33_read_write_en = (!(par_done_reg247_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg304_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg353_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg389_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg412_out | left_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_33_read_in = (!(par_done_reg228_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg286_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg338_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg379_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg406_out | top_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_23_write_out : '0;
  assign top_33_read_write_en = (!(par_done_reg228_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg286_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg338_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg379_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg406_out | top_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_33_top = (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_33_read_out : '0;
  assign pe_33_left = (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_33_read_out : '0;
  assign pe_33_go = (!pe_33_done & (!(par_done_reg270_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg324_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg368_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg399_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg418_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_32_write_in = (pe_32_done & (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_32_down : '0;
  assign down_32_write_write_en = (pe_32_done & (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_32_write_in = (pe_32_done & (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_32_right : '0;
  assign right_32_write_write_en = (pe_32_done & (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_32_read_in = (!(par_done_reg186_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg246_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg303_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg352_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg388_out | left_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_31_write_out : '0;
  assign left_32_read_write_en = (!(par_done_reg186_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg246_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg303_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg352_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg388_out | left_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_32_read_in = (!(par_done_reg168_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg227_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg285_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg337_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg378_out | top_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_22_write_out : '0;
  assign top_32_read_write_en = (!(par_done_reg168_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg227_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg285_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg337_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg378_out | top_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_32_top = (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_32_read_out : '0;
  assign pe_32_left = (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_32_read_out : '0;
  assign pe_32_go = (!pe_32_done & (!(par_done_reg210_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg269_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg323_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg367_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg398_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_31_write_in = (pe_31_done & (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_31_down : '0;
  assign down_31_write_write_en = (pe_31_done & (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_31_write_in = (pe_31_done & (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_31_right : '0;
  assign right_31_write_write_en = (pe_31_done & (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_31_read_in = (!(par_done_reg128_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg185_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg302_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg351_out | left_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_30_write_out : '0;
  assign left_31_read_write_en = (!(par_done_reg128_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg185_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg302_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg351_out | left_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_31_read_in = (!(par_done_reg113_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg226_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg284_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg336_out | top_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_21_write_out : '0;
  assign top_31_read_write_en = (!(par_done_reg113_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg226_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg284_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg336_out | top_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_31_top = (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_31_read_out : '0;
  assign pe_31_left = (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_31_read_out : '0;
  assign pe_31_go = (!pe_31_done & (!(par_done_reg151_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg268_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg322_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg366_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_30_write_in = (pe_30_done & (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_30_down : '0;
  assign down_30_write_write_en = (pe_30_done & (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_30_write_in = (pe_30_done & (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_30_right : '0;
  assign right_30_write_write_en = (pe_30_done & (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_30_read_in = (!(par_done_reg79_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg301_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? l3_read_data : '0;
  assign left_30_read_write_en = (!(par_done_reg79_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg301_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_30_read_in = (!(par_done_reg69_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg112_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg225_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg283_out | top_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_20_write_out : '0;
  assign top_30_read_write_en = (!(par_done_reg69_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg112_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg225_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg283_out | top_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_30_top = (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_30_read_out : '0;
  assign pe_30_left = (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_30_read_out : '0;
  assign pe_30_go = (!pe_30_done & (!(par_done_reg99_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg267_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg321_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_24_write_in = (pe_24_done & (!(par_done_reg266_out | down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg320_out | down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg365_out | down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg397_out | down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg417_out | down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_24_down : '0;
  assign down_24_write_write_en = (pe_24_done & (!(par_done_reg266_out | down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg320_out | down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg365_out | down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg397_out | down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg417_out | down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_24_read_in = (!(par_done_reg243_out | left_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg300_out | left_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg350_out | left_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg387_out | left_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg411_out | left_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_23_write_out : '0;
  assign left_24_read_write_en = (!(par_done_reg243_out | left_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg300_out | left_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg350_out | left_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg387_out | left_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg411_out | left_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_24_read_in = (!(par_done_reg224_out | top_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg282_out | top_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg335_out | top_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg377_out | top_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg405_out | top_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_14_write_out : '0;
  assign top_24_read_write_en = (!(par_done_reg224_out | top_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg282_out | top_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg335_out | top_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg377_out | top_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg405_out | top_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_24_top = (!(par_done_reg266_out | down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg320_out | down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg365_out | down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg397_out | down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg417_out | down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_24_read_out : '0;
  assign pe_24_left = (!(par_done_reg266_out | down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg320_out | down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg365_out | down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg397_out | down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg417_out | down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_24_read_out : '0;
  assign pe_24_go = (!pe_24_done & (!(par_done_reg266_out | down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg320_out | down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg365_out | down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg397_out | down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg417_out | down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_23_write_in = (pe_23_done & (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_23_down : '0;
  assign down_23_write_write_en = (pe_23_done & (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_23_write_in = (pe_23_done & (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_23_right : '0;
  assign right_23_write_write_en = (pe_23_done & (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_23_read_in = (!(par_done_reg183_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg242_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg299_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg349_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg386_out | left_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_22_write_out : '0;
  assign left_23_read_write_en = (!(par_done_reg183_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg242_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg299_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg349_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg386_out | left_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_23_read_in = (!(par_done_reg165_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg223_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg281_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg334_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg376_out | top_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_13_write_out : '0;
  assign top_23_read_write_en = (!(par_done_reg165_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg223_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg281_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg334_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg376_out | top_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_23_top = (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_23_read_out : '0;
  assign pe_23_left = (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_23_read_out : '0;
  assign pe_23_go = (!pe_23_done & (!(par_done_reg207_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg265_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg319_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg364_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg396_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_22_write_in = (pe_22_done & (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_22_down : '0;
  assign down_22_write_write_en = (pe_22_done & (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_22_write_in = (pe_22_done & (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_22_right : '0;
  assign right_22_write_write_en = (pe_22_done & (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_22_read_in = (!(par_done_reg126_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg182_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg298_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg348_out | left_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_21_write_out : '0;
  assign left_22_read_write_en = (!(par_done_reg126_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg182_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg298_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg348_out | left_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_22_read_in = (!(par_done_reg111_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg164_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg222_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg280_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg333_out | top_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_12_write_out : '0;
  assign top_22_read_write_en = (!(par_done_reg111_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg164_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg222_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg280_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg333_out | top_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_22_top = (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_22_read_out : '0;
  assign pe_22_left = (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_22_read_out : '0;
  assign pe_22_go = (!pe_22_done & (!(par_done_reg149_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg264_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg318_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg363_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_21_write_in = (pe_21_done & (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_21_down : '0;
  assign down_21_write_write_en = (pe_21_done & (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_21_write_in = (pe_21_done & (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_21_right : '0;
  assign right_21_write_write_en = (pe_21_done & (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_21_read_in = (!(par_done_reg78_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg125_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg181_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg297_out | left_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_20_write_out : '0;
  assign left_21_read_write_en = (!(par_done_reg78_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg125_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg181_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg297_out | left_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_21_read_in = (!(par_done_reg68_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg110_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg221_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg279_out | top_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_11_write_out : '0;
  assign top_21_read_write_en = (!(par_done_reg68_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg110_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg221_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg279_out | top_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_21_top = (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_21_read_out : '0;
  assign pe_21_left = (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_21_read_out : '0;
  assign pe_21_go = (!pe_21_done & (!(par_done_reg98_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg263_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg317_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_20_write_in = (pe_20_done & (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_20_down : '0;
  assign down_20_write_write_en = (pe_20_done & (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_20_write_in = (pe_20_done & (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_20_right : '0;
  assign right_20_write_write_en = (pe_20_done & (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_20_read_in = (!(par_done_reg45_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg180_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg239_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? l2_read_data : '0;
  assign left_20_read_write_en = (!(par_done_reg45_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg180_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg239_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_20_read_in = (!(par_done_reg39_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg162_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg220_out | top_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_10_write_out : '0;
  assign top_20_read_write_en = (!(par_done_reg39_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg162_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg220_out | top_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_20_top = (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_20_read_out : '0;
  assign pe_20_left = (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_20_read_out : '0;
  assign pe_20_go = (!pe_20_done & (!(par_done_reg59_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg262_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_14_write_in = (pe_14_done & (!(par_done_reg203_out | down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg261_out | down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg316_out | down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg362_out | down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg395_out | down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_14_down : '0;
  assign down_14_write_write_en = (pe_14_done & (!(par_done_reg203_out | down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg261_out | down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg316_out | down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg362_out | down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg395_out | down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_14_read_in = (!(par_done_reg179_out | left_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg238_out | left_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg296_out | left_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg347_out | left_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg385_out | left_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_13_write_out : '0;
  assign left_14_read_write_en = (!(par_done_reg179_out | left_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg238_out | left_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg296_out | left_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg347_out | left_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg385_out | left_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_14_read_in = (!(par_done_reg161_out | top_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg219_out | top_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg278_out | top_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg332_out | top_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg375_out | top_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_04_write_out : '0;
  assign top_14_read_write_en = (!(par_done_reg161_out | top_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg219_out | top_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg278_out | top_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg332_out | top_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg375_out | top_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_14_top = (!(par_done_reg203_out | down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg261_out | down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg316_out | down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg362_out | down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg395_out | down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_14_read_out : '0;
  assign pe_14_left = (!(par_done_reg203_out | down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg261_out | down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg316_out | down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg362_out | down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg395_out | down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_14_read_out : '0;
  assign pe_14_go = (!pe_14_done & (!(par_done_reg203_out | down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg261_out | down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg316_out | down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg362_out | down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg395_out | down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_13_write_in = (pe_13_done & (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_13_down : '0;
  assign down_13_write_write_en = (pe_13_done & (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_13_write_in = (pe_13_done & (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_13_right : '0;
  assign right_13_write_write_en = (pe_13_done & (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_13_read_in = (!(par_done_reg123_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg178_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg237_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg295_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg346_out | left_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_12_write_out : '0;
  assign left_13_read_write_en = (!(par_done_reg123_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg178_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg237_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg295_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg346_out | left_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_13_read_in = (!(par_done_reg108_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg160_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg218_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg277_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg331_out | top_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_03_write_out : '0;
  assign top_13_read_write_en = (!(par_done_reg108_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg160_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg218_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg277_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg331_out | top_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_13_top = (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_13_read_out : '0;
  assign pe_13_left = (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_13_read_out : '0;
  assign pe_13_go = (!pe_13_done & (!(par_done_reg146_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg260_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg315_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg361_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_12_write_in = (pe_12_done & (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_12_down : '0;
  assign down_12_write_write_en = (pe_12_done & (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_12_write_in = (pe_12_done & (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_12_right : '0;
  assign right_12_write_write_en = (pe_12_done & (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_12_read_in = (!(par_done_reg76_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg177_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg236_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg294_out | left_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_11_write_out : '0;
  assign left_12_read_write_en = (!(par_done_reg76_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg177_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg236_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg294_out | left_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_12_read_in = (!(par_done_reg66_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg159_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg217_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg276_out | top_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_02_write_out : '0;
  assign top_12_read_write_en = (!(par_done_reg66_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg159_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg217_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg276_out | top_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_12_top = (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_12_read_out : '0;
  assign pe_12_left = (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_12_read_out : '0;
  assign pe_12_go = (!pe_12_done & (!(par_done_reg96_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg259_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg314_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_11_write_in = (pe_11_done & (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_11_down : '0;
  assign down_11_write_write_en = (pe_11_done & (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_11_write_in = (pe_11_done & (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_11_right : '0;
  assign right_11_write_write_en = (pe_11_done & (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_11_read_in = (!(par_done_reg44_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg75_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg121_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg176_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg235_out | left_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_10_write_out : '0;
  assign left_11_read_write_en = (!(par_done_reg44_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg75_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg121_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg176_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg235_out | left_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_11_read_in = (!(par_done_reg38_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg65_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg158_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg216_out | top_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_01_write_out : '0;
  assign top_11_read_write_en = (!(par_done_reg38_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg65_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg158_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg216_out | top_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_11_top = (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_11_read_out : '0;
  assign pe_11_left = (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_11_read_out : '0;
  assign pe_11_go = (!pe_11_done & (!(par_done_reg58_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg95_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg200_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg258_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_10_write_in = (pe_10_done & (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_10_down : '0;
  assign down_10_write_write_en = (pe_10_done & (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_10_write_in = (pe_10_done & (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_10_right : '0;
  assign right_10_write_write_en = (pe_10_done & (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_10_read_in = (!(par_done_reg24_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg74_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg120_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? l1_read_data : '0;
  assign left_10_read_write_en = (!(par_done_reg24_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg74_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg120_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_10_read_in = (!(par_done_reg21_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg105_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg157_out | top_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? down_00_write_out : '0;
  assign top_10_read_write_en = (!(par_done_reg21_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg105_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg157_out | top_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_10_top = (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_10_read_out : '0;
  assign pe_10_left = (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_10_read_out : '0;
  assign pe_10_go = (!pe_10_done & (!(par_done_reg33_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg199_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign down_04_write_in = (pe_04_done & (!(par_done_reg142_out | down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg198_out | down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg257_out | down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg313_out | down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg360_out | down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_04_down : '0;
  assign down_04_write_write_en = (pe_04_done & (!(par_done_reg142_out | down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg198_out | down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg257_out | down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg313_out | down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg360_out | down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_04_read_in = (!(par_done_reg119_out | left_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg174_out | left_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg234_out | left_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg293_out | left_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg345_out | left_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_03_write_out : '0;
  assign left_04_read_write_en = (!(par_done_reg119_out | left_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg174_out | left_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg234_out | left_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg293_out | left_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg345_out | left_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_04_read_in = (!(par_done_reg104_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg156_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg215_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg275_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg330_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? t4_read_data : '0;
  assign top_04_read_write_en = (!(par_done_reg104_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg156_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg215_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg275_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg330_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_04_top = (!(par_done_reg142_out | down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg198_out | down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg257_out | down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg313_out | down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg360_out | down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_04_read_out : '0;
  assign pe_04_left = (!(par_done_reg142_out | down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg198_out | down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg257_out | down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg313_out | down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg360_out | down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_04_read_out : '0;
  assign pe_04_go = (!pe_04_done & (!(par_done_reg142_out | down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg198_out | down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg257_out | down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg313_out | down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg360_out | down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_03_write_in = (pe_03_done & (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_03_down : '0;
  assign down_03_write_write_en = (pe_03_done & (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_03_write_in = (pe_03_done & (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_03_right : '0;
  assign right_03_write_write_en = (pe_03_done & (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_03_read_in = (!(par_done_reg73_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg118_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg173_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg233_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg292_out | left_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_02_write_out : '0;
  assign left_03_read_write_en = (!(par_done_reg73_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg118_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg173_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg233_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg292_out | left_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_03_read_in = (!(par_done_reg63_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg103_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg155_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg214_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg274_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? t3_read_data : '0;
  assign top_03_read_write_en = (!(par_done_reg63_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg103_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg155_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg214_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg274_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_03_top = (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_03_read_out : '0;
  assign pe_03_left = (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_03_read_out : '0;
  assign pe_03_go = (!pe_03_done & (!(par_done_reg93_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg197_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg256_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg312_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_02_write_in = (pe_02_done & (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_02_down : '0;
  assign down_02_write_write_en = (pe_02_done & (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_02_write_in = (pe_02_done & (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_02_right : '0;
  assign right_02_write_write_en = (pe_02_done & (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_02_read_in = (!(par_done_reg42_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg117_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg172_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg232_out | left_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_01_write_out : '0;
  assign left_02_read_write_en = (!(par_done_reg42_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg117_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg172_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg232_out | left_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_02_read_in = (!(par_done_reg36_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg154_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg213_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? t2_read_data : '0;
  assign top_02_read_write_en = (!(par_done_reg36_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg154_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg213_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_02_top = (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_02_read_out : '0;
  assign pe_02_left = (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_02_read_out : '0;
  assign pe_02_go = (!pe_02_done & (!(par_done_reg56_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg196_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg255_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_01_write_in = (pe_01_done & (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_01_down : '0;
  assign down_01_write_write_en = (pe_01_done & (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_01_write_in = (pe_01_done & (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_01_right : '0;
  assign right_01_write_write_en = (pe_01_done & (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_01_read_in = (!(par_done_reg23_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg71_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg171_out | left_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? right_00_write_out : '0;
  assign left_01_read_write_en = (!(par_done_reg23_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg71_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg171_out | left_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_01_read_in = (!(par_done_reg20_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg35_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg61_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg101_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg153_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? t1_read_data : '0;
  assign top_01_read_write_en = (!(par_done_reg20_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg35_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg61_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg101_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg153_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_01_top = (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_01_read_out : '0;
  assign pe_01_left = (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_01_read_out : '0;
  assign pe_01_go = (!pe_01_done & (!(par_done_reg32_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg195_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign down_00_write_in = (pe_00_done & (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_00_down : '0;
  assign down_00_write_write_en = (pe_00_done & (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign right_00_write_in = (pe_00_done & (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_00_right : '0;
  assign right_00_write_write_en = (pe_00_done & (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign left_00_read_in = (!(par_done_reg13_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg22_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg40_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg115_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? l0_read_data : '0;
  assign left_00_read_write_en = (!(par_done_reg13_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg22_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg40_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg115_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign top_00_read_in = (!(par_done_reg12_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg19_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg34_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg100_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? t0_read_data : '0;
  assign top_00_read_write_en = (!(par_done_reg12_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg19_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg34_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg100_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign pe_00_top = (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? top_00_read_out : '0;
  assign pe_00_left = (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? left_00_read_out : '0;
  assign pe_00_go = (!pe_00_done & (!(par_done_reg18_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign l4_addr0 = (!(par_done_reg129_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg306_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg355_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? l4_idx_out : '0;
  assign l4_add_left = (!(par_done_reg89_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg194_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg254_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg311_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 3'd1 : '0;
  assign l4_add_right = (!(par_done_reg89_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg194_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg254_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg311_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? l4_idx_out : '0;
  assign l4_idx_in = (!(par_done_reg89_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg194_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg254_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg311_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? l4_add_out : (!(par_done_reg9_out | l4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l4_idx_write_en = (!(par_done_reg9_out | l4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg89_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg194_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg254_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg311_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign l3_addr0 = (!(par_done_reg79_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg301_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? l3_idx_out : '0;
  assign l3_add_left = (!(par_done_reg53_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg193_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg253_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 3'd1 : '0;
  assign l3_add_right = (!(par_done_reg53_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg193_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg253_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? l3_idx_out : '0;
  assign l3_idx_in = (!(par_done_reg53_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg193_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg253_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? l3_add_out : (!(par_done_reg8_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l3_idx_write_en = (!(par_done_reg8_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg53_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg193_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg253_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign l2_addr0 = (!(par_done_reg45_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg180_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg239_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? l2_idx_out : '0;
  assign l2_add_left = (!(par_done_reg30_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg192_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 3'd1 : '0;
  assign l2_add_right = (!(par_done_reg30_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg192_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? l2_idx_out : '0;
  assign l2_idx_in = (!(par_done_reg30_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg192_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? l2_add_out : (!(par_done_reg7_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l2_idx_write_en = (!(par_done_reg7_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg30_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg192_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign l1_addr0 = (!(par_done_reg24_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg74_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg120_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? l1_idx_out : '0;
  assign l1_add_left = (!(par_done_reg17_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 3'd1 : '0;
  assign l1_add_right = (!(par_done_reg17_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? l1_idx_out : '0;
  assign l1_idx_in = (!(par_done_reg17_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? l1_add_out : (!(par_done_reg6_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l1_idx_write_en = (!(par_done_reg6_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg17_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign l0_addr0 = (!(par_done_reg13_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg22_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg40_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg115_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? l0_idx_out : '0;
  assign l0_add_left = (!(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg15_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg26_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 3'd1 : '0;
  assign l0_add_right = (!(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg15_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg26_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? l0_idx_out : '0;
  assign l0_idx_in = (!(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg15_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg26_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? l0_add_out : (!(par_done_reg5_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l0_idx_write_en = (!(par_done_reg5_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg15_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg26_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign t4_addr0 = (!(par_done_reg104_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg156_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg215_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg275_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg330_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? t4_idx_out : '0;
  assign t4_add_left = (!(par_done_reg85_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg191_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg252_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg310_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 3'd1 : '0;
  assign t4_add_right = (!(par_done_reg85_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg191_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg252_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg310_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? t4_idx_out : '0;
  assign t4_idx_in = (!(par_done_reg85_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg191_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg252_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg310_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? t4_add_out : (!(par_done_reg4_out | t4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t4_idx_write_en = (!(par_done_reg4_out | t4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg85_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg191_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg252_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg310_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign t3_addr0 = (!(par_done_reg63_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg103_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg155_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg214_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg274_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? t3_idx_out : '0;
  assign t3_add_left = (!(par_done_reg50_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg190_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg251_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 3'd1 : '0;
  assign t3_add_right = (!(par_done_reg50_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg190_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg251_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? t3_idx_out : '0;
  assign t3_idx_in = (!(par_done_reg50_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg190_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg251_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? t3_add_out : (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t3_idx_write_en = (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg50_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg190_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg251_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign t2_addr0 = (!(par_done_reg36_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg154_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg213_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? t2_idx_out : '0;
  assign t2_add_left = (!(par_done_reg28_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg131_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg189_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 3'd1 : '0;
  assign t2_add_right = (!(par_done_reg28_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg131_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg189_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? t2_idx_out : '0;
  assign t2_idx_in = (!(par_done_reg28_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg131_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg189_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? t2_add_out : (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t2_idx_write_en = (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg28_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg131_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg189_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign t1_addr0 = (!(par_done_reg20_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg35_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg61_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg101_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg153_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? t1_idx_out : '0;
  assign t1_add_left = (!(par_done_reg16_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 3'd1 : '0;
  assign t1_add_right = (!(par_done_reg16_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? t1_idx_out : '0;
  assign t1_idx_in = (!(par_done_reg16_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? t1_add_out : (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t1_idx_write_en = (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg16_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign t0_addr0 = (!(par_done_reg12_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg19_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg34_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg100_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? t0_idx_out : '0;
  assign t0_add_left = (!(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg14_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 3'd1 : '0;
  assign t0_add_right = (!(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg14_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? t0_idx_out : '0;
  assign t0_idx_in = (!(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg14_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? t0_add_out : (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t0_idx_write_en = (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg14_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_reset0_in = par_reset0_out ? 1'd0 : (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & par_done_reg8_out & par_done_reg9_out & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_reset0_write_en = (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & par_done_reg8_out & par_done_reg9_out & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg0_in = par_reset0_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg0_write_en = (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg1_in = par_reset0_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg1_write_en = (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg2_in = par_reset0_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg2_write_en = (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg3_in = par_reset0_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg3_write_en = (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg4_in = par_reset0_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg4_write_en = (t4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg5_in = par_reset0_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg5_write_en = (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg6_in = par_reset0_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg6_write_en = (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg7_in = par_reset0_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg7_write_en = (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg8_in = par_reset0_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg8_write_en = (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg9_in = par_reset0_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg9_write_en = (l4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_reset1_in = par_reset1_out ? 1'd0 : (par_done_reg10_out & par_done_reg11_out & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_reset1_write_en = (par_done_reg10_out & par_done_reg11_out & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg10_in = par_reset1_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg10_write_en = (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg11_in = par_reset1_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg11_write_en = (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_reset2_in = par_reset2_out ? 1'd0 : (par_done_reg12_out & par_done_reg13_out & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_reset2_write_en = (par_done_reg12_out & par_done_reg13_out & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg12_in = par_reset2_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg12_write_en = (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg13_in = par_reset2_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg13_write_en = (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_reset3_in = par_reset3_out ? 1'd0 : (par_done_reg14_out & par_done_reg15_out & par_done_reg16_out & par_done_reg17_out & par_done_reg18_out & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_reset3_write_en = (par_done_reg14_out & par_done_reg15_out & par_done_reg16_out & par_done_reg17_out & par_done_reg18_out & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg14_in = par_reset3_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg14_write_en = (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg15_in = par_reset3_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg15_write_en = (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg16_in = par_reset3_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg16_write_en = (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg17_in = par_reset3_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg17_write_en = (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg18_in = par_reset3_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg18_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_reset4_in = par_reset4_out ? 1'd0 : (par_done_reg19_out & par_done_reg20_out & par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_reset4_write_en = (par_done_reg19_out & par_done_reg20_out & par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg19_in = par_reset4_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg19_write_en = (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg20_in = par_reset4_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg20_write_en = (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg21_in = par_reset4_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg21_write_en = (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg22_in = par_reset4_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg22_write_en = (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg23_in = par_reset4_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg23_write_en = (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg24_in = par_reset4_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg24_write_en = (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_reset5_in = par_reset5_out ? 1'd0 : (par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_reset5_write_en = (par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg25_in = par_reset5_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg25_write_en = (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg26_in = par_reset5_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg26_write_en = (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg27_in = par_reset5_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg27_write_en = (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg28_in = par_reset5_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg28_write_en = (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg29_in = par_reset5_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg29_write_en = (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg30_in = par_reset5_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg30_write_en = (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg31_in = par_reset5_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg31_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg32_in = par_reset5_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg32_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg33_in = par_reset5_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg33_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_reset6_in = par_reset6_out ? 1'd0 : (par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_reset6_write_en = (par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg34_in = par_reset6_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg34_write_en = (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg35_in = par_reset6_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg35_write_en = (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg36_in = par_reset6_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg36_write_en = (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg37_in = par_reset6_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg37_write_en = (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg38_in = par_reset6_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg38_write_en = (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg39_in = par_reset6_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg39_write_en = (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg40_in = par_reset6_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg40_write_en = (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg41_in = par_reset6_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg41_write_en = (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg42_in = par_reset6_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg42_write_en = (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg43_in = par_reset6_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg43_write_en = (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg44_in = par_reset6_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg44_write_en = (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg45_in = par_reset6_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg45_write_en = (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_reset7_in = par_reset7_out ? 1'd0 : (par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_reset7_write_en = (par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg46_in = par_reset7_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg46_write_en = (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg47_in = par_reset7_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg47_write_en = (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg48_in = par_reset7_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg48_write_en = (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg49_in = par_reset7_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg49_write_en = (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg50_in = par_reset7_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg50_write_en = (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg51_in = par_reset7_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg51_write_en = (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg52_in = par_reset7_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg52_write_en = (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg53_in = par_reset7_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg53_write_en = (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg54_in = par_reset7_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg54_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg55_in = par_reset7_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg55_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg56_in = par_reset7_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg56_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg57_in = par_reset7_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg57_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg58_in = par_reset7_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg58_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg59_in = par_reset7_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg59_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_reset8_in = par_reset8_out ? 1'd0 : (par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_reset8_write_en = (par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg60_in = par_reset8_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg60_write_en = (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg61_in = par_reset8_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg61_write_en = (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg62_in = par_reset8_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg62_write_en = (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg63_in = par_reset8_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg63_write_en = (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg64_in = par_reset8_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg64_write_en = (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg65_in = par_reset8_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg65_write_en = (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg66_in = par_reset8_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg66_write_en = (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg67_in = par_reset8_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg67_write_en = (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg68_in = par_reset8_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg68_write_en = (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg69_in = par_reset8_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg69_write_en = (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg70_in = par_reset8_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg70_write_en = (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg71_in = par_reset8_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg71_write_en = (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg72_in = par_reset8_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg72_write_en = (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg73_in = par_reset8_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg73_write_en = (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg74_in = par_reset8_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg74_write_en = (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg75_in = par_reset8_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg75_write_en = (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg76_in = par_reset8_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg76_write_en = (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg77_in = par_reset8_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg77_write_en = (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg78_in = par_reset8_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg78_write_en = (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg79_in = par_reset8_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg79_write_en = (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_reset9_in = par_reset9_out ? 1'd0 : (par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_reset9_write_en = (par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg80_in = par_reset9_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg80_write_en = (t0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg81_in = par_reset9_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg81_write_en = (l0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg82_in = par_reset9_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg82_write_en = (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg83_in = par_reset9_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg83_write_en = (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg84_in = par_reset9_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg84_write_en = (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg85_in = par_reset9_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg85_write_en = (t4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg86_in = par_reset9_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg86_write_en = (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg87_in = par_reset9_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg87_write_en = (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg88_in = par_reset9_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg88_write_en = (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg89_in = par_reset9_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg89_write_en = (l4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg90_in = par_reset9_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg90_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg91_in = par_reset9_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg91_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg92_in = par_reset9_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg92_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg93_in = par_reset9_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg93_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg94_in = par_reset9_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg94_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg95_in = par_reset9_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg95_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg96_in = par_reset9_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg96_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg97_in = par_reset9_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg97_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg98_in = par_reset9_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg98_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg99_in = par_reset9_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg99_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_reset10_in = par_reset10_out ? 1'd0 : (par_done_reg100_out & par_done_reg101_out & par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_reset10_write_en = (par_done_reg100_out & par_done_reg101_out & par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg100_in = par_reset10_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg100_write_en = (top_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg101_in = par_reset10_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg101_write_en = (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg102_in = par_reset10_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg102_write_en = (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg103_in = par_reset10_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg103_write_en = (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg104_in = par_reset10_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg104_write_en = (top_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg105_in = par_reset10_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg105_write_en = (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg106_in = par_reset10_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg106_write_en = (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg107_in = par_reset10_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg107_write_en = (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg108_in = par_reset10_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg108_write_en = (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg109_in = par_reset10_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg109_write_en = (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg110_in = par_reset10_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg110_write_en = (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg111_in = par_reset10_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg111_write_en = (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg112_in = par_reset10_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg112_write_en = (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg113_in = par_reset10_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg113_write_en = (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg114_in = par_reset10_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg114_write_en = (top_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg115_in = par_reset10_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg115_write_en = (left_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg116_in = par_reset10_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg116_write_en = (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg117_in = par_reset10_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg117_write_en = (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg118_in = par_reset10_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg118_write_en = (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg119_in = par_reset10_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg119_write_en = (left_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg120_in = par_reset10_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg120_write_en = (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg121_in = par_reset10_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg121_write_en = (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg122_in = par_reset10_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg122_write_en = (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg123_in = par_reset10_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg123_write_en = (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg124_in = par_reset10_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg124_write_en = (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg125_in = par_reset10_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg125_write_en = (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg126_in = par_reset10_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg126_write_en = (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg127_in = par_reset10_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg127_write_en = (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg128_in = par_reset10_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg128_write_en = (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg129_in = par_reset10_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg129_write_en = (left_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_reset11_in = par_reset11_out ? 1'd0 : (par_done_reg130_out & par_done_reg131_out & par_done_reg132_out & par_done_reg133_out & par_done_reg134_out & par_done_reg135_out & par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_reset11_write_en = (par_done_reg130_out & par_done_reg131_out & par_done_reg132_out & par_done_reg133_out & par_done_reg134_out & par_done_reg135_out & par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg130_in = par_reset11_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg130_write_en = (t1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg131_in = par_reset11_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg131_write_en = (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg132_in = par_reset11_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg132_write_en = (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg133_in = par_reset11_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg133_write_en = (t4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg134_in = par_reset11_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg134_write_en = (l1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg135_in = par_reset11_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg135_write_en = (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg136_in = par_reset11_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg136_write_en = (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg137_in = par_reset11_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg137_write_en = (l4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg138_in = par_reset11_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg138_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg139_in = par_reset11_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg139_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg140_in = par_reset11_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg140_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg141_in = par_reset11_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg141_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg142_in = par_reset11_out ? 1'd0 : (down_04_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg142_write_en = (down_04_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg143_in = par_reset11_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg143_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg144_in = par_reset11_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg144_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg145_in = par_reset11_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg145_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg146_in = par_reset11_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg146_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg147_in = par_reset11_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg147_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg148_in = par_reset11_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg148_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg149_in = par_reset11_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg149_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg150_in = par_reset11_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg150_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg151_in = par_reset11_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg151_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg152_in = par_reset11_out ? 1'd0 : (right_40_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg152_write_en = (right_40_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_reset12_in = par_reset12_out ? 1'd0 : (par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & par_done_reg158_out & par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_reset12_write_en = (par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & par_done_reg158_out & par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg153_in = par_reset12_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg153_write_en = (top_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg154_in = par_reset12_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg154_write_en = (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg155_in = par_reset12_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg155_write_en = (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg156_in = par_reset12_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg156_write_en = (top_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg157_in = par_reset12_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg157_write_en = (top_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg158_in = par_reset12_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg158_write_en = (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg159_in = par_reset12_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg159_write_en = (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg160_in = par_reset12_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg160_write_en = (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg161_in = par_reset12_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg161_write_en = (top_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg162_in = par_reset12_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg162_write_en = (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg163_in = par_reset12_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg163_write_en = (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg164_in = par_reset12_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg164_write_en = (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg165_in = par_reset12_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg165_write_en = (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg166_in = par_reset12_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg166_write_en = (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg167_in = par_reset12_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg167_write_en = (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg168_in = par_reset12_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg168_write_en = (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg169_in = par_reset12_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg169_write_en = (top_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg170_in = par_reset12_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg170_write_en = (top_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg171_in = par_reset12_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg171_write_en = (left_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg172_in = par_reset12_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg172_write_en = (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg173_in = par_reset12_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg173_write_en = (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg174_in = par_reset12_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg174_write_en = (left_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg175_in = par_reset12_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg175_write_en = (left_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg176_in = par_reset12_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg176_write_en = (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg177_in = par_reset12_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg177_write_en = (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg178_in = par_reset12_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg178_write_en = (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg179_in = par_reset12_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg179_write_en = (left_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg180_in = par_reset12_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg180_write_en = (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg181_in = par_reset12_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg181_write_en = (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg182_in = par_reset12_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg182_write_en = (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg183_in = par_reset12_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg183_write_en = (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg184_in = par_reset12_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg184_write_en = (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg185_in = par_reset12_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg185_write_en = (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg186_in = par_reset12_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg186_write_en = (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg187_in = par_reset12_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg187_write_en = (left_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg188_in = par_reset12_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg188_write_en = (left_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_reset13_in = par_reset13_out ? 1'd0 : (par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & par_done_reg201_out & par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_reset13_write_en = (par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & par_done_reg201_out & par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg189_in = par_reset13_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg189_write_en = (t2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg190_in = par_reset13_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg190_write_en = (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg191_in = par_reset13_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg191_write_en = (t4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg192_in = par_reset13_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg192_write_en = (l2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg193_in = par_reset13_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg193_write_en = (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg194_in = par_reset13_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg194_write_en = (l4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg195_in = par_reset13_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg195_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg196_in = par_reset13_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg196_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg197_in = par_reset13_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg197_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg198_in = par_reset13_out ? 1'd0 : (down_04_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg198_write_en = (down_04_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg199_in = par_reset13_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg199_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg200_in = par_reset13_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg200_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg201_in = par_reset13_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg201_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg202_in = par_reset13_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg202_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg203_in = par_reset13_out ? 1'd0 : (down_14_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg203_write_en = (down_14_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg204_in = par_reset13_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg204_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg205_in = par_reset13_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg205_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg206_in = par_reset13_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg206_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg207_in = par_reset13_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg207_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg208_in = par_reset13_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg208_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg209_in = par_reset13_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg209_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg210_in = par_reset13_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg210_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg211_in = par_reset13_out ? 1'd0 : (right_40_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg211_write_en = (right_40_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg212_in = par_reset13_out ? 1'd0 : (right_41_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg212_write_en = (right_41_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_reset14_in = par_reset14_out ? 1'd0 : (par_done_reg213_out & par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & par_done_reg229_out & par_done_reg230_out & par_done_reg231_out & par_done_reg232_out & par_done_reg233_out & par_done_reg234_out & par_done_reg235_out & par_done_reg236_out & par_done_reg237_out & par_done_reg238_out & par_done_reg239_out & par_done_reg240_out & par_done_reg241_out & par_done_reg242_out & par_done_reg243_out & par_done_reg244_out & par_done_reg245_out & par_done_reg246_out & par_done_reg247_out & par_done_reg248_out & par_done_reg249_out & par_done_reg250_out & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_reset14_write_en = (par_done_reg213_out & par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & par_done_reg229_out & par_done_reg230_out & par_done_reg231_out & par_done_reg232_out & par_done_reg233_out & par_done_reg234_out & par_done_reg235_out & par_done_reg236_out & par_done_reg237_out & par_done_reg238_out & par_done_reg239_out & par_done_reg240_out & par_done_reg241_out & par_done_reg242_out & par_done_reg243_out & par_done_reg244_out & par_done_reg245_out & par_done_reg246_out & par_done_reg247_out & par_done_reg248_out & par_done_reg249_out & par_done_reg250_out & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg213_in = par_reset14_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg213_write_en = (top_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg214_in = par_reset14_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg214_write_en = (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg215_in = par_reset14_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg215_write_en = (top_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg216_in = par_reset14_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg216_write_en = (top_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg217_in = par_reset14_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg217_write_en = (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg218_in = par_reset14_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg218_write_en = (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg219_in = par_reset14_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg219_write_en = (top_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg220_in = par_reset14_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg220_write_en = (top_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg221_in = par_reset14_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg221_write_en = (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg222_in = par_reset14_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg222_write_en = (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg223_in = par_reset14_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg223_write_en = (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg224_in = par_reset14_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg224_write_en = (top_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg225_in = par_reset14_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg225_write_en = (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg226_in = par_reset14_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg226_write_en = (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg227_in = par_reset14_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg227_write_en = (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg228_in = par_reset14_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg228_write_en = (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg229_in = par_reset14_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg229_write_en = (top_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg230_in = par_reset14_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg230_write_en = (top_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg231_in = par_reset14_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg231_write_en = (top_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg232_in = par_reset14_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg232_write_en = (left_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg233_in = par_reset14_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg233_write_en = (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg234_in = par_reset14_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg234_write_en = (left_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg235_in = par_reset14_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg235_write_en = (left_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg236_in = par_reset14_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg236_write_en = (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg237_in = par_reset14_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg237_write_en = (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg238_in = par_reset14_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg238_write_en = (left_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg239_in = par_reset14_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg239_write_en = (left_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg240_in = par_reset14_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg240_write_en = (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg241_in = par_reset14_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg241_write_en = (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg242_in = par_reset14_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg242_write_en = (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg243_in = par_reset14_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg243_write_en = (left_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg244_in = par_reset14_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg244_write_en = (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg245_in = par_reset14_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg245_write_en = (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg246_in = par_reset14_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg246_write_en = (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg247_in = par_reset14_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg247_write_en = (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg248_in = par_reset14_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg248_write_en = (left_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg249_in = par_reset14_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg249_write_en = (left_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg250_in = par_reset14_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg250_write_en = (left_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_reset15_in = par_reset15_out ? 1'd0 : (par_done_reg251_out & par_done_reg252_out & par_done_reg253_out & par_done_reg254_out & par_done_reg255_out & par_done_reg256_out & par_done_reg257_out & par_done_reg258_out & par_done_reg259_out & par_done_reg260_out & par_done_reg261_out & par_done_reg262_out & par_done_reg263_out & par_done_reg264_out & par_done_reg265_out & par_done_reg266_out & par_done_reg267_out & par_done_reg268_out & par_done_reg269_out & par_done_reg270_out & par_done_reg271_out & par_done_reg272_out & par_done_reg273_out & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_reset15_write_en = (par_done_reg251_out & par_done_reg252_out & par_done_reg253_out & par_done_reg254_out & par_done_reg255_out & par_done_reg256_out & par_done_reg257_out & par_done_reg258_out & par_done_reg259_out & par_done_reg260_out & par_done_reg261_out & par_done_reg262_out & par_done_reg263_out & par_done_reg264_out & par_done_reg265_out & par_done_reg266_out & par_done_reg267_out & par_done_reg268_out & par_done_reg269_out & par_done_reg270_out & par_done_reg271_out & par_done_reg272_out & par_done_reg273_out & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg251_in = par_reset15_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg251_write_en = (t3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg252_in = par_reset15_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg252_write_en = (t4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg253_in = par_reset15_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg253_write_en = (l3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg254_in = par_reset15_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg254_write_en = (l4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg255_in = par_reset15_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg255_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg256_in = par_reset15_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg256_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg257_in = par_reset15_out ? 1'd0 : (down_04_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg257_write_en = (down_04_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg258_in = par_reset15_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg258_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg259_in = par_reset15_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg259_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg260_in = par_reset15_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg260_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg261_in = par_reset15_out ? 1'd0 : (down_14_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg261_write_en = (down_14_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg262_in = par_reset15_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg262_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg263_in = par_reset15_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg263_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg264_in = par_reset15_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg264_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg265_in = par_reset15_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg265_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg266_in = par_reset15_out ? 1'd0 : (down_24_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg266_write_en = (down_24_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg267_in = par_reset15_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg267_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg268_in = par_reset15_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg268_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg269_in = par_reset15_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg269_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg270_in = par_reset15_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg270_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg271_in = par_reset15_out ? 1'd0 : (right_40_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg271_write_en = (right_40_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg272_in = par_reset15_out ? 1'd0 : (right_41_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg272_write_en = (right_41_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg273_in = par_reset15_out ? 1'd0 : (right_42_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg273_write_en = (right_42_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_reset16_in = par_reset16_out ? 1'd0 : (par_done_reg274_out & par_done_reg275_out & par_done_reg276_out & par_done_reg277_out & par_done_reg278_out & par_done_reg279_out & par_done_reg280_out & par_done_reg281_out & par_done_reg282_out & par_done_reg283_out & par_done_reg284_out & par_done_reg285_out & par_done_reg286_out & par_done_reg287_out & par_done_reg288_out & par_done_reg289_out & par_done_reg290_out & par_done_reg291_out & par_done_reg292_out & par_done_reg293_out & par_done_reg294_out & par_done_reg295_out & par_done_reg296_out & par_done_reg297_out & par_done_reg298_out & par_done_reg299_out & par_done_reg300_out & par_done_reg301_out & par_done_reg302_out & par_done_reg303_out & par_done_reg304_out & par_done_reg305_out & par_done_reg306_out & par_done_reg307_out & par_done_reg308_out & par_done_reg309_out & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_reset16_write_en = (par_done_reg274_out & par_done_reg275_out & par_done_reg276_out & par_done_reg277_out & par_done_reg278_out & par_done_reg279_out & par_done_reg280_out & par_done_reg281_out & par_done_reg282_out & par_done_reg283_out & par_done_reg284_out & par_done_reg285_out & par_done_reg286_out & par_done_reg287_out & par_done_reg288_out & par_done_reg289_out & par_done_reg290_out & par_done_reg291_out & par_done_reg292_out & par_done_reg293_out & par_done_reg294_out & par_done_reg295_out & par_done_reg296_out & par_done_reg297_out & par_done_reg298_out & par_done_reg299_out & par_done_reg300_out & par_done_reg301_out & par_done_reg302_out & par_done_reg303_out & par_done_reg304_out & par_done_reg305_out & par_done_reg306_out & par_done_reg307_out & par_done_reg308_out & par_done_reg309_out & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg274_in = par_reset16_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg274_write_en = (top_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg275_in = par_reset16_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg275_write_en = (top_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg276_in = par_reset16_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg276_write_en = (top_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg277_in = par_reset16_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg277_write_en = (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg278_in = par_reset16_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg278_write_en = (top_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg279_in = par_reset16_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg279_write_en = (top_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg280_in = par_reset16_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg280_write_en = (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg281_in = par_reset16_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg281_write_en = (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg282_in = par_reset16_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg282_write_en = (top_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg283_in = par_reset16_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg283_write_en = (top_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg284_in = par_reset16_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg284_write_en = (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg285_in = par_reset16_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg285_write_en = (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg286_in = par_reset16_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg286_write_en = (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg287_in = par_reset16_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg287_write_en = (top_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg288_in = par_reset16_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg288_write_en = (top_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg289_in = par_reset16_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg289_write_en = (top_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg290_in = par_reset16_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg290_write_en = (top_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg291_in = par_reset16_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg291_write_en = (top_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg292_in = par_reset16_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg292_write_en = (left_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg293_in = par_reset16_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg293_write_en = (left_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg294_in = par_reset16_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg294_write_en = (left_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg295_in = par_reset16_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg295_write_en = (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg296_in = par_reset16_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg296_write_en = (left_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg297_in = par_reset16_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg297_write_en = (left_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg298_in = par_reset16_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg298_write_en = (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg299_in = par_reset16_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg299_write_en = (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg300_in = par_reset16_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg300_write_en = (left_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg301_in = par_reset16_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg301_write_en = (left_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg302_in = par_reset16_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg302_write_en = (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg303_in = par_reset16_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg303_write_en = (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg304_in = par_reset16_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg304_write_en = (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg305_in = par_reset16_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg305_write_en = (left_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg306_in = par_reset16_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg306_write_en = (left_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg307_in = par_reset16_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg307_write_en = (left_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg308_in = par_reset16_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg308_write_en = (left_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg309_in = par_reset16_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg309_write_en = (left_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_reset17_in = par_reset17_out ? 1'd0 : (par_done_reg310_out & par_done_reg311_out & par_done_reg312_out & par_done_reg313_out & par_done_reg314_out & par_done_reg315_out & par_done_reg316_out & par_done_reg317_out & par_done_reg318_out & par_done_reg319_out & par_done_reg320_out & par_done_reg321_out & par_done_reg322_out & par_done_reg323_out & par_done_reg324_out & par_done_reg325_out & par_done_reg326_out & par_done_reg327_out & par_done_reg328_out & par_done_reg329_out & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_reset17_write_en = (par_done_reg310_out & par_done_reg311_out & par_done_reg312_out & par_done_reg313_out & par_done_reg314_out & par_done_reg315_out & par_done_reg316_out & par_done_reg317_out & par_done_reg318_out & par_done_reg319_out & par_done_reg320_out & par_done_reg321_out & par_done_reg322_out & par_done_reg323_out & par_done_reg324_out & par_done_reg325_out & par_done_reg326_out & par_done_reg327_out & par_done_reg328_out & par_done_reg329_out & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg310_in = par_reset17_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg310_write_en = (t4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg311_in = par_reset17_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg311_write_en = (l4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg312_in = par_reset17_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg312_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg313_in = par_reset17_out ? 1'd0 : (down_04_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg313_write_en = (down_04_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg314_in = par_reset17_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg314_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg315_in = par_reset17_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg315_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg316_in = par_reset17_out ? 1'd0 : (down_14_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg316_write_en = (down_14_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg317_in = par_reset17_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg317_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg318_in = par_reset17_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg318_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg319_in = par_reset17_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg319_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg320_in = par_reset17_out ? 1'd0 : (down_24_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg320_write_en = (down_24_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg321_in = par_reset17_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg321_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg322_in = par_reset17_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg322_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg323_in = par_reset17_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg323_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg324_in = par_reset17_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg324_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg325_in = par_reset17_out ? 1'd0 : (down_34_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg325_write_en = (down_34_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg326_in = par_reset17_out ? 1'd0 : (right_40_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg326_write_en = (right_40_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg327_in = par_reset17_out ? 1'd0 : (right_41_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg327_write_en = (right_41_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg328_in = par_reset17_out ? 1'd0 : (right_42_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg328_write_en = (right_42_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg329_in = par_reset17_out ? 1'd0 : (right_43_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg329_write_en = (right_43_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_reset18_in = par_reset18_out ? 1'd0 : (par_done_reg330_out & par_done_reg331_out & par_done_reg332_out & par_done_reg333_out & par_done_reg334_out & par_done_reg335_out & par_done_reg336_out & par_done_reg337_out & par_done_reg338_out & par_done_reg339_out & par_done_reg340_out & par_done_reg341_out & par_done_reg342_out & par_done_reg343_out & par_done_reg344_out & par_done_reg345_out & par_done_reg346_out & par_done_reg347_out & par_done_reg348_out & par_done_reg349_out & par_done_reg350_out & par_done_reg351_out & par_done_reg352_out & par_done_reg353_out & par_done_reg354_out & par_done_reg355_out & par_done_reg356_out & par_done_reg357_out & par_done_reg358_out & par_done_reg359_out & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_reset18_write_en = (par_done_reg330_out & par_done_reg331_out & par_done_reg332_out & par_done_reg333_out & par_done_reg334_out & par_done_reg335_out & par_done_reg336_out & par_done_reg337_out & par_done_reg338_out & par_done_reg339_out & par_done_reg340_out & par_done_reg341_out & par_done_reg342_out & par_done_reg343_out & par_done_reg344_out & par_done_reg345_out & par_done_reg346_out & par_done_reg347_out & par_done_reg348_out & par_done_reg349_out & par_done_reg350_out & par_done_reg351_out & par_done_reg352_out & par_done_reg353_out & par_done_reg354_out & par_done_reg355_out & par_done_reg356_out & par_done_reg357_out & par_done_reg358_out & par_done_reg359_out & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg330_in = par_reset18_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg330_write_en = (top_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg331_in = par_reset18_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg331_write_en = (top_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg332_in = par_reset18_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg332_write_en = (top_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg333_in = par_reset18_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg333_write_en = (top_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg334_in = par_reset18_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg334_write_en = (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg335_in = par_reset18_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg335_write_en = (top_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg336_in = par_reset18_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg336_write_en = (top_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg337_in = par_reset18_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg337_write_en = (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg338_in = par_reset18_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg338_write_en = (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg339_in = par_reset18_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg339_write_en = (top_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg340_in = par_reset18_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg340_write_en = (top_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg341_in = par_reset18_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg341_write_en = (top_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg342_in = par_reset18_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg342_write_en = (top_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg343_in = par_reset18_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg343_write_en = (top_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg344_in = par_reset18_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg344_write_en = (top_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg345_in = par_reset18_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg345_write_en = (left_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg346_in = par_reset18_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg346_write_en = (left_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg347_in = par_reset18_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg347_write_en = (left_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg348_in = par_reset18_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg348_write_en = (left_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg349_in = par_reset18_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg349_write_en = (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg350_in = par_reset18_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg350_write_en = (left_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg351_in = par_reset18_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg351_write_en = (left_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg352_in = par_reset18_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg352_write_en = (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg353_in = par_reset18_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg353_write_en = (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg354_in = par_reset18_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg354_write_en = (left_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg355_in = par_reset18_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg355_write_en = (left_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg356_in = par_reset18_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg356_write_en = (left_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg357_in = par_reset18_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg357_write_en = (left_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg358_in = par_reset18_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg358_write_en = (left_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg359_in = par_reset18_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg359_write_en = (left_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_reset19_in = par_reset19_out ? 1'd0 : (par_done_reg360_out & par_done_reg361_out & par_done_reg362_out & par_done_reg363_out & par_done_reg364_out & par_done_reg365_out & par_done_reg366_out & par_done_reg367_out & par_done_reg368_out & par_done_reg369_out & par_done_reg370_out & par_done_reg371_out & par_done_reg372_out & par_done_reg373_out & par_done_reg374_out & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_reset19_write_en = (par_done_reg360_out & par_done_reg361_out & par_done_reg362_out & par_done_reg363_out & par_done_reg364_out & par_done_reg365_out & par_done_reg366_out & par_done_reg367_out & par_done_reg368_out & par_done_reg369_out & par_done_reg370_out & par_done_reg371_out & par_done_reg372_out & par_done_reg373_out & par_done_reg374_out & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg360_in = par_reset19_out ? 1'd0 : (down_04_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg360_write_en = (down_04_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg361_in = par_reset19_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg361_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg362_in = par_reset19_out ? 1'd0 : (down_14_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg362_write_en = (down_14_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg363_in = par_reset19_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg363_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg364_in = par_reset19_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg364_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg365_in = par_reset19_out ? 1'd0 : (down_24_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg365_write_en = (down_24_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg366_in = par_reset19_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg366_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg367_in = par_reset19_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg367_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg368_in = par_reset19_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg368_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg369_in = par_reset19_out ? 1'd0 : (down_34_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg369_write_en = (down_34_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg370_in = par_reset19_out ? 1'd0 : (right_40_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg370_write_en = (right_40_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg371_in = par_reset19_out ? 1'd0 : (right_41_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg371_write_en = (right_41_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg372_in = par_reset19_out ? 1'd0 : (right_42_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg372_write_en = (right_42_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg373_in = par_reset19_out ? 1'd0 : (right_43_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg373_write_en = (right_43_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg374_in = par_reset19_out ? 1'd0 : (pe_44_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg374_write_en = (pe_44_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_reset20_in = par_reset20_out ? 1'd0 : (par_done_reg375_out & par_done_reg376_out & par_done_reg377_out & par_done_reg378_out & par_done_reg379_out & par_done_reg380_out & par_done_reg381_out & par_done_reg382_out & par_done_reg383_out & par_done_reg384_out & par_done_reg385_out & par_done_reg386_out & par_done_reg387_out & par_done_reg388_out & par_done_reg389_out & par_done_reg390_out & par_done_reg391_out & par_done_reg392_out & par_done_reg393_out & par_done_reg394_out & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_reset20_write_en = (par_done_reg375_out & par_done_reg376_out & par_done_reg377_out & par_done_reg378_out & par_done_reg379_out & par_done_reg380_out & par_done_reg381_out & par_done_reg382_out & par_done_reg383_out & par_done_reg384_out & par_done_reg385_out & par_done_reg386_out & par_done_reg387_out & par_done_reg388_out & par_done_reg389_out & par_done_reg390_out & par_done_reg391_out & par_done_reg392_out & par_done_reg393_out & par_done_reg394_out & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg375_in = par_reset20_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg375_write_en = (top_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg376_in = par_reset20_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg376_write_en = (top_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg377_in = par_reset20_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg377_write_en = (top_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg378_in = par_reset20_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg378_write_en = (top_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg379_in = par_reset20_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg379_write_en = (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg380_in = par_reset20_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg380_write_en = (top_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg381_in = par_reset20_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg381_write_en = (top_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg382_in = par_reset20_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg382_write_en = (top_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg383_in = par_reset20_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg383_write_en = (top_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg384_in = par_reset20_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg384_write_en = (top_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg385_in = par_reset20_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg385_write_en = (left_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg386_in = par_reset20_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg386_write_en = (left_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg387_in = par_reset20_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg387_write_en = (left_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg388_in = par_reset20_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg388_write_en = (left_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg389_in = par_reset20_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg389_write_en = (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg390_in = par_reset20_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg390_write_en = (left_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg391_in = par_reset20_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg391_write_en = (left_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg392_in = par_reset20_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg392_write_en = (left_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg393_in = par_reset20_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg393_write_en = (left_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg394_in = par_reset20_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg394_write_en = (left_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_reset21_in = par_reset21_out ? 1'd0 : (par_done_reg395_out & par_done_reg396_out & par_done_reg397_out & par_done_reg398_out & par_done_reg399_out & par_done_reg400_out & par_done_reg401_out & par_done_reg402_out & par_done_reg403_out & par_done_reg404_out & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_reset21_write_en = (par_done_reg395_out & par_done_reg396_out & par_done_reg397_out & par_done_reg398_out & par_done_reg399_out & par_done_reg400_out & par_done_reg401_out & par_done_reg402_out & par_done_reg403_out & par_done_reg404_out & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg395_in = par_reset21_out ? 1'd0 : (down_14_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg395_write_en = (down_14_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg396_in = par_reset21_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg396_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg397_in = par_reset21_out ? 1'd0 : (down_24_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg397_write_en = (down_24_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg398_in = par_reset21_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg398_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg399_in = par_reset21_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg399_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg400_in = par_reset21_out ? 1'd0 : (down_34_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg400_write_en = (down_34_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg401_in = par_reset21_out ? 1'd0 : (right_41_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg401_write_en = (right_41_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg402_in = par_reset21_out ? 1'd0 : (right_42_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg402_write_en = (right_42_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg403_in = par_reset21_out ? 1'd0 : (right_43_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg403_write_en = (right_43_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg404_in = par_reset21_out ? 1'd0 : (pe_44_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg404_write_en = (pe_44_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_reset22_in = par_reset22_out ? 1'd0 : (par_done_reg405_out & par_done_reg406_out & par_done_reg407_out & par_done_reg408_out & par_done_reg409_out & par_done_reg410_out & par_done_reg411_out & par_done_reg412_out & par_done_reg413_out & par_done_reg414_out & par_done_reg415_out & par_done_reg416_out & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_reset22_write_en = (par_done_reg405_out & par_done_reg406_out & par_done_reg407_out & par_done_reg408_out & par_done_reg409_out & par_done_reg410_out & par_done_reg411_out & par_done_reg412_out & par_done_reg413_out & par_done_reg414_out & par_done_reg415_out & par_done_reg416_out & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg405_in = par_reset22_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg405_write_en = (top_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg406_in = par_reset22_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg406_write_en = (top_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg407_in = par_reset22_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg407_write_en = (top_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg408_in = par_reset22_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg408_write_en = (top_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg409_in = par_reset22_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg409_write_en = (top_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg410_in = par_reset22_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg410_write_en = (top_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg411_in = par_reset22_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg411_write_en = (left_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg412_in = par_reset22_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg412_write_en = (left_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg413_in = par_reset22_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg413_write_en = (left_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg414_in = par_reset22_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg414_write_en = (left_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg415_in = par_reset22_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg415_write_en = (left_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg416_in = par_reset22_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg416_write_en = (left_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_reset23_in = par_reset23_out ? 1'd0 : (par_done_reg417_out & par_done_reg418_out & par_done_reg419_out & par_done_reg420_out & par_done_reg421_out & par_done_reg422_out & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_reset23_write_en = (par_done_reg417_out & par_done_reg418_out & par_done_reg419_out & par_done_reg420_out & par_done_reg421_out & par_done_reg422_out & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg417_in = par_reset23_out ? 1'd0 : (down_24_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg417_write_en = (down_24_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg418_in = par_reset23_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg418_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg419_in = par_reset23_out ? 1'd0 : (down_34_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg419_write_en = (down_34_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg420_in = par_reset23_out ? 1'd0 : (right_42_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg420_write_en = (right_42_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg421_in = par_reset23_out ? 1'd0 : (right_43_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg421_write_en = (right_43_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg422_in = par_reset23_out ? 1'd0 : (pe_44_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg422_write_en = (pe_44_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_reset24_in = par_reset24_out ? 1'd0 : (par_done_reg423_out & par_done_reg424_out & par_done_reg425_out & par_done_reg426_out & par_done_reg427_out & par_done_reg428_out & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_reset24_write_en = (par_done_reg423_out & par_done_reg424_out & par_done_reg425_out & par_done_reg426_out & par_done_reg427_out & par_done_reg428_out & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg423_in = par_reset24_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg423_write_en = (top_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg424_in = par_reset24_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg424_write_en = (top_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg425_in = par_reset24_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg425_write_en = (top_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg426_in = par_reset24_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg426_write_en = (left_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg427_in = par_reset24_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg427_write_en = (left_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg428_in = par_reset24_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg428_write_en = (left_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_reset25_in = par_reset25_out ? 1'd0 : (par_done_reg429_out & par_done_reg430_out & par_done_reg431_out & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_reset25_write_en = (par_done_reg429_out & par_done_reg430_out & par_done_reg431_out & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg429_in = par_reset25_out ? 1'd0 : (down_34_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg429_write_en = (down_34_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg430_in = par_reset25_out ? 1'd0 : (right_43_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg430_write_en = (right_43_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg431_in = par_reset25_out ? 1'd0 : (pe_44_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg431_write_en = (pe_44_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_reset26_in = par_reset26_out ? 1'd0 : (par_done_reg432_out & par_done_reg433_out & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_reset26_write_en = (par_done_reg432_out & par_done_reg433_out & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg432_in = par_reset26_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg432_write_en = (top_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg433_in = par_reset26_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg433_write_en = (left_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_reset27_in = par_reset27_out ? 1'd0 : (par_done_reg434_out & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_reset27_write_en = (par_done_reg434_out & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg434_in = par_reset27_out ? 1'd0 : (pe_44_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg434_write_en = (pe_44_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd0 & par_reset0_out & go) ? 32'd1 : (fsm0_out == 32'd53) ? 32'd0 : (fsm0_out == 32'd52 & out_mem_done & go) ? 32'd53 : (fsm0_out == 32'd51 & out_mem_done & go) ? 32'd52 : (fsm0_out == 32'd50 & out_mem_done & go) ? 32'd51 : (fsm0_out == 32'd49 & out_mem_done & go) ? 32'd50 : (fsm0_out == 32'd48 & out_mem_done & go) ? 32'd49 : (fsm0_out == 32'd47 & out_mem_done & go) ? 32'd48 : (fsm0_out == 32'd46 & out_mem_done & go) ? 32'd47 : (fsm0_out == 32'd45 & out_mem_done & go) ? 32'd46 : (fsm0_out == 32'd44 & out_mem_done & go) ? 32'd45 : (fsm0_out == 32'd43 & out_mem_done & go) ? 32'd44 : (fsm0_out == 32'd42 & out_mem_done & go) ? 32'd43 : (fsm0_out == 32'd41 & out_mem_done & go) ? 32'd42 : (fsm0_out == 32'd40 & out_mem_done & go) ? 32'd41 : (fsm0_out == 32'd39 & out_mem_done & go) ? 32'd40 : (fsm0_out == 32'd38 & out_mem_done & go) ? 32'd39 : (fsm0_out == 32'd37 & out_mem_done & go) ? 32'd38 : (fsm0_out == 32'd36 & out_mem_done & go) ? 32'd37 : (fsm0_out == 32'd35 & out_mem_done & go) ? 32'd36 : (fsm0_out == 32'd34 & out_mem_done & go) ? 32'd35 : (fsm0_out == 32'd33 & out_mem_done & go) ? 32'd34 : (fsm0_out == 32'd32 & out_mem_done & go) ? 32'd33 : (fsm0_out == 32'd31 & out_mem_done & go) ? 32'd32 : (fsm0_out == 32'd30 & out_mem_done & go) ? 32'd31 : (fsm0_out == 32'd29 & out_mem_done & go) ? 32'd30 : (fsm0_out == 32'd28 & out_mem_done & go) ? 32'd29 : (fsm0_out == 32'd27 & par_reset27_out & go) ? 32'd28 : (fsm0_out == 32'd26 & par_reset26_out & go) ? 32'd27 : (fsm0_out == 32'd25 & par_reset25_out & go) ? 32'd26 : (fsm0_out == 32'd24 & par_reset24_out & go) ? 32'd25 : (fsm0_out == 32'd23 & par_reset23_out & go) ? 32'd24 : (fsm0_out == 32'd22 & par_reset22_out & go) ? 32'd23 : (fsm0_out == 32'd21 & par_reset21_out & go) ? 32'd22 : (fsm0_out == 32'd20 & par_reset20_out & go) ? 32'd21 : (fsm0_out == 32'd19 & par_reset19_out & go) ? 32'd20 : (fsm0_out == 32'd18 & par_reset18_out & go) ? 32'd19 : (fsm0_out == 32'd17 & par_reset17_out & go) ? 32'd18 : (fsm0_out == 32'd16 & par_reset16_out & go) ? 32'd17 : (fsm0_out == 32'd15 & par_reset15_out & go) ? 32'd16 : (fsm0_out == 32'd14 & par_reset14_out & go) ? 32'd15 : (fsm0_out == 32'd13 & par_reset13_out & go) ? 32'd14 : (fsm0_out == 32'd12 & par_reset12_out & go) ? 32'd13 : (fsm0_out == 32'd11 & par_reset11_out & go) ? 32'd12 : (fsm0_out == 32'd10 & par_reset10_out & go) ? 32'd11 : (fsm0_out == 32'd9 & par_reset9_out & go) ? 32'd10 : (fsm0_out == 32'd8 & par_reset8_out & go) ? 32'd9 : (fsm0_out == 32'd7 & par_reset7_out & go) ? 32'd8 : (fsm0_out == 32'd6 & par_reset6_out & go) ? 32'd7 : (fsm0_out == 32'd5 & par_reset5_out & go) ? 32'd6 : (fsm0_out == 32'd4 & par_reset4_out & go) ? 32'd5 : (fsm0_out == 32'd3 & par_reset3_out & go) ? 32'd4 : (fsm0_out == 32'd2 & par_reset2_out & go) ? 32'd3 : (fsm0_out == 32'd1 & par_reset1_out & go) ? 32'd2 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & par_reset0_out & go | fsm0_out == 32'd1 & par_reset1_out & go | fsm0_out == 32'd2 & par_reset2_out & go | fsm0_out == 32'd3 & par_reset3_out & go | fsm0_out == 32'd4 & par_reset4_out & go | fsm0_out == 32'd5 & par_reset5_out & go | fsm0_out == 32'd6 & par_reset6_out & go | fsm0_out == 32'd7 & par_reset7_out & go | fsm0_out == 32'd8 & par_reset8_out & go | fsm0_out == 32'd9 & par_reset9_out & go | fsm0_out == 32'd10 & par_reset10_out & go | fsm0_out == 32'd11 & par_reset11_out & go | fsm0_out == 32'd12 & par_reset12_out & go | fsm0_out == 32'd13 & par_reset13_out & go | fsm0_out == 32'd14 & par_reset14_out & go | fsm0_out == 32'd15 & par_reset15_out & go | fsm0_out == 32'd16 & par_reset16_out & go | fsm0_out == 32'd17 & par_reset17_out & go | fsm0_out == 32'd18 & par_reset18_out & go | fsm0_out == 32'd19 & par_reset19_out & go | fsm0_out == 32'd20 & par_reset20_out & go | fsm0_out == 32'd21 & par_reset21_out & go | fsm0_out == 32'd22 & par_reset22_out & go | fsm0_out == 32'd23 & par_reset23_out & go | fsm0_out == 32'd24 & par_reset24_out & go | fsm0_out == 32'd25 & par_reset25_out & go | fsm0_out == 32'd26 & par_reset26_out & go | fsm0_out == 32'd27 & par_reset27_out & go | fsm0_out == 32'd28 & out_mem_done & go | fsm0_out == 32'd29 & out_mem_done & go | fsm0_out == 32'd30 & out_mem_done & go | fsm0_out == 32'd31 & out_mem_done & go | fsm0_out == 32'd32 & out_mem_done & go | fsm0_out == 32'd33 & out_mem_done & go | fsm0_out == 32'd34 & out_mem_done & go | fsm0_out == 32'd35 & out_mem_done & go | fsm0_out == 32'd36 & out_mem_done & go | fsm0_out == 32'd37 & out_mem_done & go | fsm0_out == 32'd38 & out_mem_done & go | fsm0_out == 32'd39 & out_mem_done & go | fsm0_out == 32'd40 & out_mem_done & go | fsm0_out == 32'd41 & out_mem_done & go | fsm0_out == 32'd42 & out_mem_done & go | fsm0_out == 32'd43 & out_mem_done & go | fsm0_out == 32'd44 & out_mem_done & go | fsm0_out == 32'd45 & out_mem_done & go | fsm0_out == 32'd46 & out_mem_done & go | fsm0_out == 32'd47 & out_mem_done & go | fsm0_out == 32'd48 & out_mem_done & go | fsm0_out == 32'd49 & out_mem_done & go | fsm0_out == 32'd50 & out_mem_done & go | fsm0_out == 32'd51 & out_mem_done & go | fsm0_out == 32'd52 & out_mem_done & go | fsm0_out == 32'd53) ? 1'd1 : '0;
endmodule // end main