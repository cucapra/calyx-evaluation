/* verilator lint_off WIDTH */
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule

module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule

module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

// Component Signature
module mac_pe (
      input wire [31:0] top,
      input wire [31:0] left,
      input wire go,
      input wire clk,
      output wire [31:0] down,
      output wire [31:0] right,
      output wire [31:0] out,
      output wire done
  );
  
  // Structure wire declarations
  wire [31:0] mul_left;
  wire [31:0] mul_right;
  wire mul_go;
  wire mul_clk;
  wire [31:0] mul_out;
  wire mul_done;
  wire [31:0] add_left;
  wire [31:0] add_right;
  wire [31:0] add_out;
  wire [31:0] mul_reg_in;
  wire mul_reg_write_en;
  wire mul_reg_clk;
  wire [31:0] mul_reg_out;
  wire mul_reg_done;
  wire [31:0] acc_in;
  wire acc_write_en;
  wire acc_clk;
  wire [31:0] acc_out;
  wire acc_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_mult_pipe #(32) mul (
      .left(mul_left),
      .right(mul_right),
      .go(mul_go),
      .clk(clk),
      .out(mul_out),
      .done(mul_done)
  );
  
  std_add #(32) add (
      .left(add_left),
      .right(add_right),
      .out(add_out)
  );
  
  std_reg #(32) mul_reg (
      .in(mul_reg_in),
      .write_en(mul_reg_write_en),
      .clk(clk),
      .out(mul_reg_out),
      .done(mul_reg_done)
  );
  
  std_reg #(32) acc (
      .in(acc_in),
      .write_en(acc_write_en),
      .clk(clk),
      .out(acc_out),
      .done(acc_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign down = top;
  assign right = left;
  assign out = acc_out;
  assign done = (fsm0_out == 32'd2) ? 1'd1 : '0;
  assign mul_left = (fsm0_out == 32'd0 & !mul_reg_done & go) ? top : '0;
  assign mul_right = (fsm0_out == 32'd0 & !mul_reg_done & go) ? left : '0;
  assign mul_go = (!mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign add_left = (fsm0_out == 32'd1 & !acc_done & go) ? acc_out : '0;
  assign add_right = (fsm0_out == 32'd1 & !acc_done & go) ? mul_reg_out : '0;
  assign mul_reg_in = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? mul_out : '0;
  assign mul_reg_write_en = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign acc_in = (fsm0_out == 32'd1 & !acc_done & go) ? add_out : '0;
  assign acc_write_en = (fsm0_out == 32'd1 & !acc_done & go) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd1 & acc_done & go) ? 32'd2 : (fsm0_out == 32'd0 & mul_reg_done & go) ? 32'd1 : (fsm0_out == 32'd2) ? 32'd0 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & mul_reg_done & go | fsm0_out == 32'd1 & acc_done & go | fsm0_out == 32'd2) ? 1'd1 : '0;
endmodule // end mac_pe
// Component Signature
module main (
      input wire go,
      input wire clk,
      input wire [31:0] out_mem_read_data,
      input wire out_mem_done,
      output wire done,
      output wire [1:0] out_mem_addr0,
      output wire [1:0] out_mem_addr1,
      output wire [31:0] out_mem_write_data,
      output wire out_mem_write_en
  );
  
  // Structure wire declarations
  wire [31:0] left_22_read_in;
  wire left_22_read_write_en;
  wire left_22_read_clk;
  wire [31:0] left_22_read_out;
  wire left_22_read_done;
  wire [31:0] top_22_read_in;
  wire top_22_read_write_en;
  wire top_22_read_clk;
  wire [31:0] top_22_read_out;
  wire top_22_read_done;
  wire [31:0] pe_22_top;
  wire [31:0] pe_22_left;
  wire pe_22_go;
  wire pe_22_clk;
  wire [31:0] pe_22_down;
  wire [31:0] pe_22_right;
  wire [31:0] pe_22_out;
  wire pe_22_done;
  wire [31:0] right_21_write_in;
  wire right_21_write_write_en;
  wire right_21_write_clk;
  wire [31:0] right_21_write_out;
  wire right_21_write_done;
  wire [31:0] left_21_read_in;
  wire left_21_read_write_en;
  wire left_21_read_clk;
  wire [31:0] left_21_read_out;
  wire left_21_read_done;
  wire [31:0] top_21_read_in;
  wire top_21_read_write_en;
  wire top_21_read_clk;
  wire [31:0] top_21_read_out;
  wire top_21_read_done;
  wire [31:0] pe_21_top;
  wire [31:0] pe_21_left;
  wire pe_21_go;
  wire pe_21_clk;
  wire [31:0] pe_21_down;
  wire [31:0] pe_21_right;
  wire [31:0] pe_21_out;
  wire pe_21_done;
  wire [31:0] right_20_write_in;
  wire right_20_write_write_en;
  wire right_20_write_clk;
  wire [31:0] right_20_write_out;
  wire right_20_write_done;
  wire [31:0] left_20_read_in;
  wire left_20_read_write_en;
  wire left_20_read_clk;
  wire [31:0] left_20_read_out;
  wire left_20_read_done;
  wire [31:0] top_20_read_in;
  wire top_20_read_write_en;
  wire top_20_read_clk;
  wire [31:0] top_20_read_out;
  wire top_20_read_done;
  wire [31:0] pe_20_top;
  wire [31:0] pe_20_left;
  wire pe_20_go;
  wire pe_20_clk;
  wire [31:0] pe_20_down;
  wire [31:0] pe_20_right;
  wire [31:0] pe_20_out;
  wire pe_20_done;
  wire [31:0] down_12_write_in;
  wire down_12_write_write_en;
  wire down_12_write_clk;
  wire [31:0] down_12_write_out;
  wire down_12_write_done;
  wire [31:0] left_12_read_in;
  wire left_12_read_write_en;
  wire left_12_read_clk;
  wire [31:0] left_12_read_out;
  wire left_12_read_done;
  wire [31:0] top_12_read_in;
  wire top_12_read_write_en;
  wire top_12_read_clk;
  wire [31:0] top_12_read_out;
  wire top_12_read_done;
  wire [31:0] pe_12_top;
  wire [31:0] pe_12_left;
  wire pe_12_go;
  wire pe_12_clk;
  wire [31:0] pe_12_down;
  wire [31:0] pe_12_right;
  wire [31:0] pe_12_out;
  wire pe_12_done;
  wire [31:0] down_11_write_in;
  wire down_11_write_write_en;
  wire down_11_write_clk;
  wire [31:0] down_11_write_out;
  wire down_11_write_done;
  wire [31:0] right_11_write_in;
  wire right_11_write_write_en;
  wire right_11_write_clk;
  wire [31:0] right_11_write_out;
  wire right_11_write_done;
  wire [31:0] left_11_read_in;
  wire left_11_read_write_en;
  wire left_11_read_clk;
  wire [31:0] left_11_read_out;
  wire left_11_read_done;
  wire [31:0] top_11_read_in;
  wire top_11_read_write_en;
  wire top_11_read_clk;
  wire [31:0] top_11_read_out;
  wire top_11_read_done;
  wire [31:0] pe_11_top;
  wire [31:0] pe_11_left;
  wire pe_11_go;
  wire pe_11_clk;
  wire [31:0] pe_11_down;
  wire [31:0] pe_11_right;
  wire [31:0] pe_11_out;
  wire pe_11_done;
  wire [31:0] down_10_write_in;
  wire down_10_write_write_en;
  wire down_10_write_clk;
  wire [31:0] down_10_write_out;
  wire down_10_write_done;
  wire [31:0] right_10_write_in;
  wire right_10_write_write_en;
  wire right_10_write_clk;
  wire [31:0] right_10_write_out;
  wire right_10_write_done;
  wire [31:0] left_10_read_in;
  wire left_10_read_write_en;
  wire left_10_read_clk;
  wire [31:0] left_10_read_out;
  wire left_10_read_done;
  wire [31:0] top_10_read_in;
  wire top_10_read_write_en;
  wire top_10_read_clk;
  wire [31:0] top_10_read_out;
  wire top_10_read_done;
  wire [31:0] pe_10_top;
  wire [31:0] pe_10_left;
  wire pe_10_go;
  wire pe_10_clk;
  wire [31:0] pe_10_down;
  wire [31:0] pe_10_right;
  wire [31:0] pe_10_out;
  wire pe_10_done;
  wire [31:0] down_02_write_in;
  wire down_02_write_write_en;
  wire down_02_write_clk;
  wire [31:0] down_02_write_out;
  wire down_02_write_done;
  wire [31:0] left_02_read_in;
  wire left_02_read_write_en;
  wire left_02_read_clk;
  wire [31:0] left_02_read_out;
  wire left_02_read_done;
  wire [31:0] top_02_read_in;
  wire top_02_read_write_en;
  wire top_02_read_clk;
  wire [31:0] top_02_read_out;
  wire top_02_read_done;
  wire [31:0] pe_02_top;
  wire [31:0] pe_02_left;
  wire pe_02_go;
  wire pe_02_clk;
  wire [31:0] pe_02_down;
  wire [31:0] pe_02_right;
  wire [31:0] pe_02_out;
  wire pe_02_done;
  wire [31:0] down_01_write_in;
  wire down_01_write_write_en;
  wire down_01_write_clk;
  wire [31:0] down_01_write_out;
  wire down_01_write_done;
  wire [31:0] right_01_write_in;
  wire right_01_write_write_en;
  wire right_01_write_clk;
  wire [31:0] right_01_write_out;
  wire right_01_write_done;
  wire [31:0] left_01_read_in;
  wire left_01_read_write_en;
  wire left_01_read_clk;
  wire [31:0] left_01_read_out;
  wire left_01_read_done;
  wire [31:0] top_01_read_in;
  wire top_01_read_write_en;
  wire top_01_read_clk;
  wire [31:0] top_01_read_out;
  wire top_01_read_done;
  wire [31:0] pe_01_top;
  wire [31:0] pe_01_left;
  wire pe_01_go;
  wire pe_01_clk;
  wire [31:0] pe_01_down;
  wire [31:0] pe_01_right;
  wire [31:0] pe_01_out;
  wire pe_01_done;
  wire [31:0] down_00_write_in;
  wire down_00_write_write_en;
  wire down_00_write_clk;
  wire [31:0] down_00_write_out;
  wire down_00_write_done;
  wire [31:0] right_00_write_in;
  wire right_00_write_write_en;
  wire right_00_write_clk;
  wire [31:0] right_00_write_out;
  wire right_00_write_done;
  wire [31:0] left_00_read_in;
  wire left_00_read_write_en;
  wire left_00_read_clk;
  wire [31:0] left_00_read_out;
  wire left_00_read_done;
  wire [31:0] top_00_read_in;
  wire top_00_read_write_en;
  wire top_00_read_clk;
  wire [31:0] top_00_read_out;
  wire top_00_read_done;
  wire [31:0] pe_00_top;
  wire [31:0] pe_00_left;
  wire pe_00_go;
  wire pe_00_clk;
  wire [31:0] pe_00_down;
  wire [31:0] pe_00_right;
  wire [31:0] pe_00_out;
  wire pe_00_done;
  wire [1:0] l2_addr0;
  wire [31:0] l2_write_data;
  wire l2_write_en;
  wire l2_clk;
  wire [31:0] l2_read_data;
  wire l2_done;
  wire [1:0] l2_add_left;
  wire [1:0] l2_add_right;
  wire [1:0] l2_add_out;
  wire [1:0] l2_idx_in;
  wire l2_idx_write_en;
  wire l2_idx_clk;
  wire [1:0] l2_idx_out;
  wire l2_idx_done;
  wire [1:0] l1_addr0;
  wire [31:0] l1_write_data;
  wire l1_write_en;
  wire l1_clk;
  wire [31:0] l1_read_data;
  wire l1_done;
  wire [1:0] l1_add_left;
  wire [1:0] l1_add_right;
  wire [1:0] l1_add_out;
  wire [1:0] l1_idx_in;
  wire l1_idx_write_en;
  wire l1_idx_clk;
  wire [1:0] l1_idx_out;
  wire l1_idx_done;
  wire [1:0] l0_addr0;
  wire [31:0] l0_write_data;
  wire l0_write_en;
  wire l0_clk;
  wire [31:0] l0_read_data;
  wire l0_done;
  wire [1:0] l0_add_left;
  wire [1:0] l0_add_right;
  wire [1:0] l0_add_out;
  wire [1:0] l0_idx_in;
  wire l0_idx_write_en;
  wire l0_idx_clk;
  wire [1:0] l0_idx_out;
  wire l0_idx_done;
  wire [1:0] t2_addr0;
  wire [31:0] t2_write_data;
  wire t2_write_en;
  wire t2_clk;
  wire [31:0] t2_read_data;
  wire t2_done;
  wire [1:0] t2_add_left;
  wire [1:0] t2_add_right;
  wire [1:0] t2_add_out;
  wire [1:0] t2_idx_in;
  wire t2_idx_write_en;
  wire t2_idx_clk;
  wire [1:0] t2_idx_out;
  wire t2_idx_done;
  wire [1:0] t1_addr0;
  wire [31:0] t1_write_data;
  wire t1_write_en;
  wire t1_clk;
  wire [31:0] t1_read_data;
  wire t1_done;
  wire [1:0] t1_add_left;
  wire [1:0] t1_add_right;
  wire [1:0] t1_add_out;
  wire [1:0] t1_idx_in;
  wire t1_idx_write_en;
  wire t1_idx_clk;
  wire [1:0] t1_idx_out;
  wire t1_idx_done;
  wire [1:0] t0_addr0;
  wire [31:0] t0_write_data;
  wire t0_write_en;
  wire t0_clk;
  wire [31:0] t0_read_data;
  wire t0_done;
  wire [1:0] t0_add_left;
  wire [1:0] t0_add_right;
  wire [1:0] t0_add_out;
  wire [1:0] t0_idx_in;
  wire t0_idx_write_en;
  wire t0_idx_clk;
  wire [1:0] t0_idx_out;
  wire t0_idx_done;
  wire par_reset0_in;
  wire par_reset0_write_en;
  wire par_reset0_clk;
  wire par_reset0_out;
  wire par_reset0_done;
  wire par_done_reg0_in;
  wire par_done_reg0_write_en;
  wire par_done_reg0_clk;
  wire par_done_reg0_out;
  wire par_done_reg0_done;
  wire par_done_reg1_in;
  wire par_done_reg1_write_en;
  wire par_done_reg1_clk;
  wire par_done_reg1_out;
  wire par_done_reg1_done;
  wire par_done_reg2_in;
  wire par_done_reg2_write_en;
  wire par_done_reg2_clk;
  wire par_done_reg2_out;
  wire par_done_reg2_done;
  wire par_done_reg3_in;
  wire par_done_reg3_write_en;
  wire par_done_reg3_clk;
  wire par_done_reg3_out;
  wire par_done_reg3_done;
  wire par_done_reg4_in;
  wire par_done_reg4_write_en;
  wire par_done_reg4_clk;
  wire par_done_reg4_out;
  wire par_done_reg4_done;
  wire par_done_reg5_in;
  wire par_done_reg5_write_en;
  wire par_done_reg5_clk;
  wire par_done_reg5_out;
  wire par_done_reg5_done;
  wire par_reset1_in;
  wire par_reset1_write_en;
  wire par_reset1_clk;
  wire par_reset1_out;
  wire par_reset1_done;
  wire par_done_reg6_in;
  wire par_done_reg6_write_en;
  wire par_done_reg6_clk;
  wire par_done_reg6_out;
  wire par_done_reg6_done;
  wire par_done_reg7_in;
  wire par_done_reg7_write_en;
  wire par_done_reg7_clk;
  wire par_done_reg7_out;
  wire par_done_reg7_done;
  wire par_reset2_in;
  wire par_reset2_write_en;
  wire par_reset2_clk;
  wire par_reset2_out;
  wire par_reset2_done;
  wire par_done_reg8_in;
  wire par_done_reg8_write_en;
  wire par_done_reg8_clk;
  wire par_done_reg8_out;
  wire par_done_reg8_done;
  wire par_done_reg9_in;
  wire par_done_reg9_write_en;
  wire par_done_reg9_clk;
  wire par_done_reg9_out;
  wire par_done_reg9_done;
  wire par_reset3_in;
  wire par_reset3_write_en;
  wire par_reset3_clk;
  wire par_reset3_out;
  wire par_reset3_done;
  wire par_done_reg10_in;
  wire par_done_reg10_write_en;
  wire par_done_reg10_clk;
  wire par_done_reg10_out;
  wire par_done_reg10_done;
  wire par_done_reg11_in;
  wire par_done_reg11_write_en;
  wire par_done_reg11_clk;
  wire par_done_reg11_out;
  wire par_done_reg11_done;
  wire par_done_reg12_in;
  wire par_done_reg12_write_en;
  wire par_done_reg12_clk;
  wire par_done_reg12_out;
  wire par_done_reg12_done;
  wire par_done_reg13_in;
  wire par_done_reg13_write_en;
  wire par_done_reg13_clk;
  wire par_done_reg13_out;
  wire par_done_reg13_done;
  wire par_done_reg14_in;
  wire par_done_reg14_write_en;
  wire par_done_reg14_clk;
  wire par_done_reg14_out;
  wire par_done_reg14_done;
  wire par_reset4_in;
  wire par_reset4_write_en;
  wire par_reset4_clk;
  wire par_reset4_out;
  wire par_reset4_done;
  wire par_done_reg15_in;
  wire par_done_reg15_write_en;
  wire par_done_reg15_clk;
  wire par_done_reg15_out;
  wire par_done_reg15_done;
  wire par_done_reg16_in;
  wire par_done_reg16_write_en;
  wire par_done_reg16_clk;
  wire par_done_reg16_out;
  wire par_done_reg16_done;
  wire par_done_reg17_in;
  wire par_done_reg17_write_en;
  wire par_done_reg17_clk;
  wire par_done_reg17_out;
  wire par_done_reg17_done;
  wire par_done_reg18_in;
  wire par_done_reg18_write_en;
  wire par_done_reg18_clk;
  wire par_done_reg18_out;
  wire par_done_reg18_done;
  wire par_done_reg19_in;
  wire par_done_reg19_write_en;
  wire par_done_reg19_clk;
  wire par_done_reg19_out;
  wire par_done_reg19_done;
  wire par_done_reg20_in;
  wire par_done_reg20_write_en;
  wire par_done_reg20_clk;
  wire par_done_reg20_out;
  wire par_done_reg20_done;
  wire par_reset5_in;
  wire par_reset5_write_en;
  wire par_reset5_clk;
  wire par_reset5_out;
  wire par_reset5_done;
  wire par_done_reg21_in;
  wire par_done_reg21_write_en;
  wire par_done_reg21_clk;
  wire par_done_reg21_out;
  wire par_done_reg21_done;
  wire par_done_reg22_in;
  wire par_done_reg22_write_en;
  wire par_done_reg22_clk;
  wire par_done_reg22_out;
  wire par_done_reg22_done;
  wire par_done_reg23_in;
  wire par_done_reg23_write_en;
  wire par_done_reg23_clk;
  wire par_done_reg23_out;
  wire par_done_reg23_done;
  wire par_done_reg24_in;
  wire par_done_reg24_write_en;
  wire par_done_reg24_clk;
  wire par_done_reg24_out;
  wire par_done_reg24_done;
  wire par_done_reg25_in;
  wire par_done_reg25_write_en;
  wire par_done_reg25_clk;
  wire par_done_reg25_out;
  wire par_done_reg25_done;
  wire par_done_reg26_in;
  wire par_done_reg26_write_en;
  wire par_done_reg26_clk;
  wire par_done_reg26_out;
  wire par_done_reg26_done;
  wire par_done_reg27_in;
  wire par_done_reg27_write_en;
  wire par_done_reg27_clk;
  wire par_done_reg27_out;
  wire par_done_reg27_done;
  wire par_done_reg28_in;
  wire par_done_reg28_write_en;
  wire par_done_reg28_clk;
  wire par_done_reg28_out;
  wire par_done_reg28_done;
  wire par_done_reg29_in;
  wire par_done_reg29_write_en;
  wire par_done_reg29_clk;
  wire par_done_reg29_out;
  wire par_done_reg29_done;
  wire par_reset6_in;
  wire par_reset6_write_en;
  wire par_reset6_clk;
  wire par_reset6_out;
  wire par_reset6_done;
  wire par_done_reg30_in;
  wire par_done_reg30_write_en;
  wire par_done_reg30_clk;
  wire par_done_reg30_out;
  wire par_done_reg30_done;
  wire par_done_reg31_in;
  wire par_done_reg31_write_en;
  wire par_done_reg31_clk;
  wire par_done_reg31_out;
  wire par_done_reg31_done;
  wire par_done_reg32_in;
  wire par_done_reg32_write_en;
  wire par_done_reg32_clk;
  wire par_done_reg32_out;
  wire par_done_reg32_done;
  wire par_done_reg33_in;
  wire par_done_reg33_write_en;
  wire par_done_reg33_clk;
  wire par_done_reg33_out;
  wire par_done_reg33_done;
  wire par_done_reg34_in;
  wire par_done_reg34_write_en;
  wire par_done_reg34_clk;
  wire par_done_reg34_out;
  wire par_done_reg34_done;
  wire par_done_reg35_in;
  wire par_done_reg35_write_en;
  wire par_done_reg35_clk;
  wire par_done_reg35_out;
  wire par_done_reg35_done;
  wire par_done_reg36_in;
  wire par_done_reg36_write_en;
  wire par_done_reg36_clk;
  wire par_done_reg36_out;
  wire par_done_reg36_done;
  wire par_done_reg37_in;
  wire par_done_reg37_write_en;
  wire par_done_reg37_clk;
  wire par_done_reg37_out;
  wire par_done_reg37_done;
  wire par_done_reg38_in;
  wire par_done_reg38_write_en;
  wire par_done_reg38_clk;
  wire par_done_reg38_out;
  wire par_done_reg38_done;
  wire par_done_reg39_in;
  wire par_done_reg39_write_en;
  wire par_done_reg39_clk;
  wire par_done_reg39_out;
  wire par_done_reg39_done;
  wire par_done_reg40_in;
  wire par_done_reg40_write_en;
  wire par_done_reg40_clk;
  wire par_done_reg40_out;
  wire par_done_reg40_done;
  wire par_done_reg41_in;
  wire par_done_reg41_write_en;
  wire par_done_reg41_clk;
  wire par_done_reg41_out;
  wire par_done_reg41_done;
  wire par_reset7_in;
  wire par_reset7_write_en;
  wire par_reset7_clk;
  wire par_reset7_out;
  wire par_reset7_done;
  wire par_done_reg42_in;
  wire par_done_reg42_write_en;
  wire par_done_reg42_clk;
  wire par_done_reg42_out;
  wire par_done_reg42_done;
  wire par_done_reg43_in;
  wire par_done_reg43_write_en;
  wire par_done_reg43_clk;
  wire par_done_reg43_out;
  wire par_done_reg43_done;
  wire par_done_reg44_in;
  wire par_done_reg44_write_en;
  wire par_done_reg44_clk;
  wire par_done_reg44_out;
  wire par_done_reg44_done;
  wire par_done_reg45_in;
  wire par_done_reg45_write_en;
  wire par_done_reg45_clk;
  wire par_done_reg45_out;
  wire par_done_reg45_done;
  wire par_done_reg46_in;
  wire par_done_reg46_write_en;
  wire par_done_reg46_clk;
  wire par_done_reg46_out;
  wire par_done_reg46_done;
  wire par_done_reg47_in;
  wire par_done_reg47_write_en;
  wire par_done_reg47_clk;
  wire par_done_reg47_out;
  wire par_done_reg47_done;
  wire par_done_reg48_in;
  wire par_done_reg48_write_en;
  wire par_done_reg48_clk;
  wire par_done_reg48_out;
  wire par_done_reg48_done;
  wire par_done_reg49_in;
  wire par_done_reg49_write_en;
  wire par_done_reg49_clk;
  wire par_done_reg49_out;
  wire par_done_reg49_done;
  wire par_done_reg50_in;
  wire par_done_reg50_write_en;
  wire par_done_reg50_clk;
  wire par_done_reg50_out;
  wire par_done_reg50_done;
  wire par_done_reg51_in;
  wire par_done_reg51_write_en;
  wire par_done_reg51_clk;
  wire par_done_reg51_out;
  wire par_done_reg51_done;
  wire par_reset8_in;
  wire par_reset8_write_en;
  wire par_reset8_clk;
  wire par_reset8_out;
  wire par_reset8_done;
  wire par_done_reg52_in;
  wire par_done_reg52_write_en;
  wire par_done_reg52_clk;
  wire par_done_reg52_out;
  wire par_done_reg52_done;
  wire par_done_reg53_in;
  wire par_done_reg53_write_en;
  wire par_done_reg53_clk;
  wire par_done_reg53_out;
  wire par_done_reg53_done;
  wire par_done_reg54_in;
  wire par_done_reg54_write_en;
  wire par_done_reg54_clk;
  wire par_done_reg54_out;
  wire par_done_reg54_done;
  wire par_done_reg55_in;
  wire par_done_reg55_write_en;
  wire par_done_reg55_clk;
  wire par_done_reg55_out;
  wire par_done_reg55_done;
  wire par_done_reg56_in;
  wire par_done_reg56_write_en;
  wire par_done_reg56_clk;
  wire par_done_reg56_out;
  wire par_done_reg56_done;
  wire par_done_reg57_in;
  wire par_done_reg57_write_en;
  wire par_done_reg57_clk;
  wire par_done_reg57_out;
  wire par_done_reg57_done;
  wire par_done_reg58_in;
  wire par_done_reg58_write_en;
  wire par_done_reg58_clk;
  wire par_done_reg58_out;
  wire par_done_reg58_done;
  wire par_done_reg59_in;
  wire par_done_reg59_write_en;
  wire par_done_reg59_clk;
  wire par_done_reg59_out;
  wire par_done_reg59_done;
  wire par_done_reg60_in;
  wire par_done_reg60_write_en;
  wire par_done_reg60_clk;
  wire par_done_reg60_out;
  wire par_done_reg60_done;
  wire par_done_reg61_in;
  wire par_done_reg61_write_en;
  wire par_done_reg61_clk;
  wire par_done_reg61_out;
  wire par_done_reg61_done;
  wire par_done_reg62_in;
  wire par_done_reg62_write_en;
  wire par_done_reg62_clk;
  wire par_done_reg62_out;
  wire par_done_reg62_done;
  wire par_done_reg63_in;
  wire par_done_reg63_write_en;
  wire par_done_reg63_clk;
  wire par_done_reg63_out;
  wire par_done_reg63_done;
  wire par_done_reg64_in;
  wire par_done_reg64_write_en;
  wire par_done_reg64_clk;
  wire par_done_reg64_out;
  wire par_done_reg64_done;
  wire par_done_reg65_in;
  wire par_done_reg65_write_en;
  wire par_done_reg65_clk;
  wire par_done_reg65_out;
  wire par_done_reg65_done;
  wire par_reset9_in;
  wire par_reset9_write_en;
  wire par_reset9_clk;
  wire par_reset9_out;
  wire par_reset9_done;
  wire par_done_reg66_in;
  wire par_done_reg66_write_en;
  wire par_done_reg66_clk;
  wire par_done_reg66_out;
  wire par_done_reg66_done;
  wire par_done_reg67_in;
  wire par_done_reg67_write_en;
  wire par_done_reg67_clk;
  wire par_done_reg67_out;
  wire par_done_reg67_done;
  wire par_done_reg68_in;
  wire par_done_reg68_write_en;
  wire par_done_reg68_clk;
  wire par_done_reg68_out;
  wire par_done_reg68_done;
  wire par_done_reg69_in;
  wire par_done_reg69_write_en;
  wire par_done_reg69_clk;
  wire par_done_reg69_out;
  wire par_done_reg69_done;
  wire par_done_reg70_in;
  wire par_done_reg70_write_en;
  wire par_done_reg70_clk;
  wire par_done_reg70_out;
  wire par_done_reg70_done;
  wire par_done_reg71_in;
  wire par_done_reg71_write_en;
  wire par_done_reg71_clk;
  wire par_done_reg71_out;
  wire par_done_reg71_done;
  wire par_done_reg72_in;
  wire par_done_reg72_write_en;
  wire par_done_reg72_clk;
  wire par_done_reg72_out;
  wire par_done_reg72_done;
  wire par_done_reg73_in;
  wire par_done_reg73_write_en;
  wire par_done_reg73_clk;
  wire par_done_reg73_out;
  wire par_done_reg73_done;
  wire par_done_reg74_in;
  wire par_done_reg74_write_en;
  wire par_done_reg74_clk;
  wire par_done_reg74_out;
  wire par_done_reg74_done;
  wire par_reset10_in;
  wire par_reset10_write_en;
  wire par_reset10_clk;
  wire par_reset10_out;
  wire par_reset10_done;
  wire par_done_reg75_in;
  wire par_done_reg75_write_en;
  wire par_done_reg75_clk;
  wire par_done_reg75_out;
  wire par_done_reg75_done;
  wire par_done_reg76_in;
  wire par_done_reg76_write_en;
  wire par_done_reg76_clk;
  wire par_done_reg76_out;
  wire par_done_reg76_done;
  wire par_done_reg77_in;
  wire par_done_reg77_write_en;
  wire par_done_reg77_clk;
  wire par_done_reg77_out;
  wire par_done_reg77_done;
  wire par_done_reg78_in;
  wire par_done_reg78_write_en;
  wire par_done_reg78_clk;
  wire par_done_reg78_out;
  wire par_done_reg78_done;
  wire par_done_reg79_in;
  wire par_done_reg79_write_en;
  wire par_done_reg79_clk;
  wire par_done_reg79_out;
  wire par_done_reg79_done;
  wire par_done_reg80_in;
  wire par_done_reg80_write_en;
  wire par_done_reg80_clk;
  wire par_done_reg80_out;
  wire par_done_reg80_done;
  wire par_done_reg81_in;
  wire par_done_reg81_write_en;
  wire par_done_reg81_clk;
  wire par_done_reg81_out;
  wire par_done_reg81_done;
  wire par_done_reg82_in;
  wire par_done_reg82_write_en;
  wire par_done_reg82_clk;
  wire par_done_reg82_out;
  wire par_done_reg82_done;
  wire par_done_reg83_in;
  wire par_done_reg83_write_en;
  wire par_done_reg83_clk;
  wire par_done_reg83_out;
  wire par_done_reg83_done;
  wire par_done_reg84_in;
  wire par_done_reg84_write_en;
  wire par_done_reg84_clk;
  wire par_done_reg84_out;
  wire par_done_reg84_done;
  wire par_done_reg85_in;
  wire par_done_reg85_write_en;
  wire par_done_reg85_clk;
  wire par_done_reg85_out;
  wire par_done_reg85_done;
  wire par_done_reg86_in;
  wire par_done_reg86_write_en;
  wire par_done_reg86_clk;
  wire par_done_reg86_out;
  wire par_done_reg86_done;
  wire par_reset11_in;
  wire par_reset11_write_en;
  wire par_reset11_clk;
  wire par_reset11_out;
  wire par_reset11_done;
  wire par_done_reg87_in;
  wire par_done_reg87_write_en;
  wire par_done_reg87_clk;
  wire par_done_reg87_out;
  wire par_done_reg87_done;
  wire par_done_reg88_in;
  wire par_done_reg88_write_en;
  wire par_done_reg88_clk;
  wire par_done_reg88_out;
  wire par_done_reg88_done;
  wire par_done_reg89_in;
  wire par_done_reg89_write_en;
  wire par_done_reg89_clk;
  wire par_done_reg89_out;
  wire par_done_reg89_done;
  wire par_done_reg90_in;
  wire par_done_reg90_write_en;
  wire par_done_reg90_clk;
  wire par_done_reg90_out;
  wire par_done_reg90_done;
  wire par_done_reg91_in;
  wire par_done_reg91_write_en;
  wire par_done_reg91_clk;
  wire par_done_reg91_out;
  wire par_done_reg91_done;
  wire par_done_reg92_in;
  wire par_done_reg92_write_en;
  wire par_done_reg92_clk;
  wire par_done_reg92_out;
  wire par_done_reg92_done;
  wire par_reset12_in;
  wire par_reset12_write_en;
  wire par_reset12_clk;
  wire par_reset12_out;
  wire par_reset12_done;
  wire par_done_reg93_in;
  wire par_done_reg93_write_en;
  wire par_done_reg93_clk;
  wire par_done_reg93_out;
  wire par_done_reg93_done;
  wire par_done_reg94_in;
  wire par_done_reg94_write_en;
  wire par_done_reg94_clk;
  wire par_done_reg94_out;
  wire par_done_reg94_done;
  wire par_done_reg95_in;
  wire par_done_reg95_write_en;
  wire par_done_reg95_clk;
  wire par_done_reg95_out;
  wire par_done_reg95_done;
  wire par_done_reg96_in;
  wire par_done_reg96_write_en;
  wire par_done_reg96_clk;
  wire par_done_reg96_out;
  wire par_done_reg96_done;
  wire par_done_reg97_in;
  wire par_done_reg97_write_en;
  wire par_done_reg97_clk;
  wire par_done_reg97_out;
  wire par_done_reg97_done;
  wire par_done_reg98_in;
  wire par_done_reg98_write_en;
  wire par_done_reg98_clk;
  wire par_done_reg98_out;
  wire par_done_reg98_done;
  wire par_reset13_in;
  wire par_reset13_write_en;
  wire par_reset13_clk;
  wire par_reset13_out;
  wire par_reset13_done;
  wire par_done_reg99_in;
  wire par_done_reg99_write_en;
  wire par_done_reg99_clk;
  wire par_done_reg99_out;
  wire par_done_reg99_done;
  wire par_done_reg100_in;
  wire par_done_reg100_write_en;
  wire par_done_reg100_clk;
  wire par_done_reg100_out;
  wire par_done_reg100_done;
  wire par_done_reg101_in;
  wire par_done_reg101_write_en;
  wire par_done_reg101_clk;
  wire par_done_reg101_out;
  wire par_done_reg101_done;
  wire par_reset14_in;
  wire par_reset14_write_en;
  wire par_reset14_clk;
  wire par_reset14_out;
  wire par_reset14_done;
  wire par_done_reg102_in;
  wire par_done_reg102_write_en;
  wire par_done_reg102_clk;
  wire par_done_reg102_out;
  wire par_done_reg102_done;
  wire par_done_reg103_in;
  wire par_done_reg103_write_en;
  wire par_done_reg103_clk;
  wire par_done_reg103_out;
  wire par_done_reg103_done;
  wire par_reset15_in;
  wire par_reset15_write_en;
  wire par_reset15_clk;
  wire par_reset15_out;
  wire par_reset15_done;
  wire par_done_reg104_in;
  wire par_done_reg104_write_en;
  wire par_done_reg104_clk;
  wire par_done_reg104_out;
  wire par_done_reg104_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_reg #(32) left_22_read (
      .in(left_22_read_in),
      .write_en(left_22_read_write_en),
      .clk(clk),
      .out(left_22_read_out),
      .done(left_22_read_done)
  );
  
  std_reg #(32) top_22_read (
      .in(top_22_read_in),
      .write_en(top_22_read_write_en),
      .clk(clk),
      .out(top_22_read_out),
      .done(top_22_read_done)
  );
  
  mac_pe #() pe_22 (
      .top(pe_22_top),
      .left(pe_22_left),
      .go(pe_22_go),
      .clk(clk),
      .down(pe_22_down),
      .right(pe_22_right),
      .out(pe_22_out),
      .done(pe_22_done)
  );
  
  std_reg #(32) right_21_write (
      .in(right_21_write_in),
      .write_en(right_21_write_write_en),
      .clk(clk),
      .out(right_21_write_out),
      .done(right_21_write_done)
  );
  
  std_reg #(32) left_21_read (
      .in(left_21_read_in),
      .write_en(left_21_read_write_en),
      .clk(clk),
      .out(left_21_read_out),
      .done(left_21_read_done)
  );
  
  std_reg #(32) top_21_read (
      .in(top_21_read_in),
      .write_en(top_21_read_write_en),
      .clk(clk),
      .out(top_21_read_out),
      .done(top_21_read_done)
  );
  
  mac_pe #() pe_21 (
      .top(pe_21_top),
      .left(pe_21_left),
      .go(pe_21_go),
      .clk(clk),
      .down(pe_21_down),
      .right(pe_21_right),
      .out(pe_21_out),
      .done(pe_21_done)
  );
  
  std_reg #(32) right_20_write (
      .in(right_20_write_in),
      .write_en(right_20_write_write_en),
      .clk(clk),
      .out(right_20_write_out),
      .done(right_20_write_done)
  );
  
  std_reg #(32) left_20_read (
      .in(left_20_read_in),
      .write_en(left_20_read_write_en),
      .clk(clk),
      .out(left_20_read_out),
      .done(left_20_read_done)
  );
  
  std_reg #(32) top_20_read (
      .in(top_20_read_in),
      .write_en(top_20_read_write_en),
      .clk(clk),
      .out(top_20_read_out),
      .done(top_20_read_done)
  );
  
  mac_pe #() pe_20 (
      .top(pe_20_top),
      .left(pe_20_left),
      .go(pe_20_go),
      .clk(clk),
      .down(pe_20_down),
      .right(pe_20_right),
      .out(pe_20_out),
      .done(pe_20_done)
  );
  
  std_reg #(32) down_12_write (
      .in(down_12_write_in),
      .write_en(down_12_write_write_en),
      .clk(clk),
      .out(down_12_write_out),
      .done(down_12_write_done)
  );
  
  std_reg #(32) left_12_read (
      .in(left_12_read_in),
      .write_en(left_12_read_write_en),
      .clk(clk),
      .out(left_12_read_out),
      .done(left_12_read_done)
  );
  
  std_reg #(32) top_12_read (
      .in(top_12_read_in),
      .write_en(top_12_read_write_en),
      .clk(clk),
      .out(top_12_read_out),
      .done(top_12_read_done)
  );
  
  mac_pe #() pe_12 (
      .top(pe_12_top),
      .left(pe_12_left),
      .go(pe_12_go),
      .clk(clk),
      .down(pe_12_down),
      .right(pe_12_right),
      .out(pe_12_out),
      .done(pe_12_done)
  );
  
  std_reg #(32) down_11_write (
      .in(down_11_write_in),
      .write_en(down_11_write_write_en),
      .clk(clk),
      .out(down_11_write_out),
      .done(down_11_write_done)
  );
  
  std_reg #(32) right_11_write (
      .in(right_11_write_in),
      .write_en(right_11_write_write_en),
      .clk(clk),
      .out(right_11_write_out),
      .done(right_11_write_done)
  );
  
  std_reg #(32) left_11_read (
      .in(left_11_read_in),
      .write_en(left_11_read_write_en),
      .clk(clk),
      .out(left_11_read_out),
      .done(left_11_read_done)
  );
  
  std_reg #(32) top_11_read (
      .in(top_11_read_in),
      .write_en(top_11_read_write_en),
      .clk(clk),
      .out(top_11_read_out),
      .done(top_11_read_done)
  );
  
  mac_pe #() pe_11 (
      .top(pe_11_top),
      .left(pe_11_left),
      .go(pe_11_go),
      .clk(clk),
      .down(pe_11_down),
      .right(pe_11_right),
      .out(pe_11_out),
      .done(pe_11_done)
  );
  
  std_reg #(32) down_10_write (
      .in(down_10_write_in),
      .write_en(down_10_write_write_en),
      .clk(clk),
      .out(down_10_write_out),
      .done(down_10_write_done)
  );
  
  std_reg #(32) right_10_write (
      .in(right_10_write_in),
      .write_en(right_10_write_write_en),
      .clk(clk),
      .out(right_10_write_out),
      .done(right_10_write_done)
  );
  
  std_reg #(32) left_10_read (
      .in(left_10_read_in),
      .write_en(left_10_read_write_en),
      .clk(clk),
      .out(left_10_read_out),
      .done(left_10_read_done)
  );
  
  std_reg #(32) top_10_read (
      .in(top_10_read_in),
      .write_en(top_10_read_write_en),
      .clk(clk),
      .out(top_10_read_out),
      .done(top_10_read_done)
  );
  
  mac_pe #() pe_10 (
      .top(pe_10_top),
      .left(pe_10_left),
      .go(pe_10_go),
      .clk(clk),
      .down(pe_10_down),
      .right(pe_10_right),
      .out(pe_10_out),
      .done(pe_10_done)
  );
  
  std_reg #(32) down_02_write (
      .in(down_02_write_in),
      .write_en(down_02_write_write_en),
      .clk(clk),
      .out(down_02_write_out),
      .done(down_02_write_done)
  );
  
  std_reg #(32) left_02_read (
      .in(left_02_read_in),
      .write_en(left_02_read_write_en),
      .clk(clk),
      .out(left_02_read_out),
      .done(left_02_read_done)
  );
  
  std_reg #(32) top_02_read (
      .in(top_02_read_in),
      .write_en(top_02_read_write_en),
      .clk(clk),
      .out(top_02_read_out),
      .done(top_02_read_done)
  );
  
  mac_pe #() pe_02 (
      .top(pe_02_top),
      .left(pe_02_left),
      .go(pe_02_go),
      .clk(clk),
      .down(pe_02_down),
      .right(pe_02_right),
      .out(pe_02_out),
      .done(pe_02_done)
  );
  
  std_reg #(32) down_01_write (
      .in(down_01_write_in),
      .write_en(down_01_write_write_en),
      .clk(clk),
      .out(down_01_write_out),
      .done(down_01_write_done)
  );
  
  std_reg #(32) right_01_write (
      .in(right_01_write_in),
      .write_en(right_01_write_write_en),
      .clk(clk),
      .out(right_01_write_out),
      .done(right_01_write_done)
  );
  
  std_reg #(32) left_01_read (
      .in(left_01_read_in),
      .write_en(left_01_read_write_en),
      .clk(clk),
      .out(left_01_read_out),
      .done(left_01_read_done)
  );
  
  std_reg #(32) top_01_read (
      .in(top_01_read_in),
      .write_en(top_01_read_write_en),
      .clk(clk),
      .out(top_01_read_out),
      .done(top_01_read_done)
  );
  
  mac_pe #() pe_01 (
      .top(pe_01_top),
      .left(pe_01_left),
      .go(pe_01_go),
      .clk(clk),
      .down(pe_01_down),
      .right(pe_01_right),
      .out(pe_01_out),
      .done(pe_01_done)
  );
  
  std_reg #(32) down_00_write (
      .in(down_00_write_in),
      .write_en(down_00_write_write_en),
      .clk(clk),
      .out(down_00_write_out),
      .done(down_00_write_done)
  );
  
  std_reg #(32) right_00_write (
      .in(right_00_write_in),
      .write_en(right_00_write_write_en),
      .clk(clk),
      .out(right_00_write_out),
      .done(right_00_write_done)
  );
  
  std_reg #(32) left_00_read (
      .in(left_00_read_in),
      .write_en(left_00_read_write_en),
      .clk(clk),
      .out(left_00_read_out),
      .done(left_00_read_done)
  );
  
  std_reg #(32) top_00_read (
      .in(top_00_read_in),
      .write_en(top_00_read_write_en),
      .clk(clk),
      .out(top_00_read_out),
      .done(top_00_read_done)
  );
  
  mac_pe #() pe_00 (
      .top(pe_00_top),
      .left(pe_00_left),
      .go(pe_00_go),
      .clk(clk),
      .down(pe_00_down),
      .right(pe_00_right),
      .out(pe_00_out),
      .done(pe_00_done)
  );
  
  std_mem_d1 #(32, 3, 2) l2 (
      .addr0(l2_addr0),
      .write_data(l2_write_data),
      .write_en(l2_write_en),
      .clk(clk),
      .read_data(l2_read_data),
      .done(l2_done)
  );
  
  std_add #(2) l2_add (
      .left(l2_add_left),
      .right(l2_add_right),
      .out(l2_add_out)
  );
  
  std_reg #(2) l2_idx (
      .in(l2_idx_in),
      .write_en(l2_idx_write_en),
      .clk(clk),
      .out(l2_idx_out),
      .done(l2_idx_done)
  );
  
  std_mem_d1 #(32, 3, 2) l1 (
      .addr0(l1_addr0),
      .write_data(l1_write_data),
      .write_en(l1_write_en),
      .clk(clk),
      .read_data(l1_read_data),
      .done(l1_done)
  );
  
  std_add #(2) l1_add (
      .left(l1_add_left),
      .right(l1_add_right),
      .out(l1_add_out)
  );
  
  std_reg #(2) l1_idx (
      .in(l1_idx_in),
      .write_en(l1_idx_write_en),
      .clk(clk),
      .out(l1_idx_out),
      .done(l1_idx_done)
  );
  
  std_mem_d1 #(32, 3, 2) l0 (
      .addr0(l0_addr0),
      .write_data(l0_write_data),
      .write_en(l0_write_en),
      .clk(clk),
      .read_data(l0_read_data),
      .done(l0_done)
  );
  
  std_add #(2) l0_add (
      .left(l0_add_left),
      .right(l0_add_right),
      .out(l0_add_out)
  );
  
  std_reg #(2) l0_idx (
      .in(l0_idx_in),
      .write_en(l0_idx_write_en),
      .clk(clk),
      .out(l0_idx_out),
      .done(l0_idx_done)
  );
  
  std_mem_d1 #(32, 3, 2) t2 (
      .addr0(t2_addr0),
      .write_data(t2_write_data),
      .write_en(t2_write_en),
      .clk(clk),
      .read_data(t2_read_data),
      .done(t2_done)
  );
  
  std_add #(2) t2_add (
      .left(t2_add_left),
      .right(t2_add_right),
      .out(t2_add_out)
  );
  
  std_reg #(2) t2_idx (
      .in(t2_idx_in),
      .write_en(t2_idx_write_en),
      .clk(clk),
      .out(t2_idx_out),
      .done(t2_idx_done)
  );
  
  std_mem_d1 #(32, 3, 2) t1 (
      .addr0(t1_addr0),
      .write_data(t1_write_data),
      .write_en(t1_write_en),
      .clk(clk),
      .read_data(t1_read_data),
      .done(t1_done)
  );
  
  std_add #(2) t1_add (
      .left(t1_add_left),
      .right(t1_add_right),
      .out(t1_add_out)
  );
  
  std_reg #(2) t1_idx (
      .in(t1_idx_in),
      .write_en(t1_idx_write_en),
      .clk(clk),
      .out(t1_idx_out),
      .done(t1_idx_done)
  );
  
  std_mem_d1 #(32, 3, 2) t0 (
      .addr0(t0_addr0),
      .write_data(t0_write_data),
      .write_en(t0_write_en),
      .clk(clk),
      .read_data(t0_read_data),
      .done(t0_done)
  );
  
  std_add #(2) t0_add (
      .left(t0_add_left),
      .right(t0_add_right),
      .out(t0_add_out)
  );
  
  std_reg #(2) t0_idx (
      .in(t0_idx_in),
      .write_en(t0_idx_write_en),
      .clk(clk),
      .out(t0_idx_out),
      .done(t0_idx_done)
  );
  
  std_reg #(1) par_reset0 (
      .in(par_reset0_in),
      .write_en(par_reset0_write_en),
      .clk(clk),
      .out(par_reset0_out),
      .done(par_reset0_done)
  );
  
  std_reg #(1) par_done_reg0 (
      .in(par_done_reg0_in),
      .write_en(par_done_reg0_write_en),
      .clk(clk),
      .out(par_done_reg0_out),
      .done(par_done_reg0_done)
  );
  
  std_reg #(1) par_done_reg1 (
      .in(par_done_reg1_in),
      .write_en(par_done_reg1_write_en),
      .clk(clk),
      .out(par_done_reg1_out),
      .done(par_done_reg1_done)
  );
  
  std_reg #(1) par_done_reg2 (
      .in(par_done_reg2_in),
      .write_en(par_done_reg2_write_en),
      .clk(clk),
      .out(par_done_reg2_out),
      .done(par_done_reg2_done)
  );
  
  std_reg #(1) par_done_reg3 (
      .in(par_done_reg3_in),
      .write_en(par_done_reg3_write_en),
      .clk(clk),
      .out(par_done_reg3_out),
      .done(par_done_reg3_done)
  );
  
  std_reg #(1) par_done_reg4 (
      .in(par_done_reg4_in),
      .write_en(par_done_reg4_write_en),
      .clk(clk),
      .out(par_done_reg4_out),
      .done(par_done_reg4_done)
  );
  
  std_reg #(1) par_done_reg5 (
      .in(par_done_reg5_in),
      .write_en(par_done_reg5_write_en),
      .clk(clk),
      .out(par_done_reg5_out),
      .done(par_done_reg5_done)
  );
  
  std_reg #(1) par_reset1 (
      .in(par_reset1_in),
      .write_en(par_reset1_write_en),
      .clk(clk),
      .out(par_reset1_out),
      .done(par_reset1_done)
  );
  
  std_reg #(1) par_done_reg6 (
      .in(par_done_reg6_in),
      .write_en(par_done_reg6_write_en),
      .clk(clk),
      .out(par_done_reg6_out),
      .done(par_done_reg6_done)
  );
  
  std_reg #(1) par_done_reg7 (
      .in(par_done_reg7_in),
      .write_en(par_done_reg7_write_en),
      .clk(clk),
      .out(par_done_reg7_out),
      .done(par_done_reg7_done)
  );
  
  std_reg #(1) par_reset2 (
      .in(par_reset2_in),
      .write_en(par_reset2_write_en),
      .clk(clk),
      .out(par_reset2_out),
      .done(par_reset2_done)
  );
  
  std_reg #(1) par_done_reg8 (
      .in(par_done_reg8_in),
      .write_en(par_done_reg8_write_en),
      .clk(clk),
      .out(par_done_reg8_out),
      .done(par_done_reg8_done)
  );
  
  std_reg #(1) par_done_reg9 (
      .in(par_done_reg9_in),
      .write_en(par_done_reg9_write_en),
      .clk(clk),
      .out(par_done_reg9_out),
      .done(par_done_reg9_done)
  );
  
  std_reg #(1) par_reset3 (
      .in(par_reset3_in),
      .write_en(par_reset3_write_en),
      .clk(clk),
      .out(par_reset3_out),
      .done(par_reset3_done)
  );
  
  std_reg #(1) par_done_reg10 (
      .in(par_done_reg10_in),
      .write_en(par_done_reg10_write_en),
      .clk(clk),
      .out(par_done_reg10_out),
      .done(par_done_reg10_done)
  );
  
  std_reg #(1) par_done_reg11 (
      .in(par_done_reg11_in),
      .write_en(par_done_reg11_write_en),
      .clk(clk),
      .out(par_done_reg11_out),
      .done(par_done_reg11_done)
  );
  
  std_reg #(1) par_done_reg12 (
      .in(par_done_reg12_in),
      .write_en(par_done_reg12_write_en),
      .clk(clk),
      .out(par_done_reg12_out),
      .done(par_done_reg12_done)
  );
  
  std_reg #(1) par_done_reg13 (
      .in(par_done_reg13_in),
      .write_en(par_done_reg13_write_en),
      .clk(clk),
      .out(par_done_reg13_out),
      .done(par_done_reg13_done)
  );
  
  std_reg #(1) par_done_reg14 (
      .in(par_done_reg14_in),
      .write_en(par_done_reg14_write_en),
      .clk(clk),
      .out(par_done_reg14_out),
      .done(par_done_reg14_done)
  );
  
  std_reg #(1) par_reset4 (
      .in(par_reset4_in),
      .write_en(par_reset4_write_en),
      .clk(clk),
      .out(par_reset4_out),
      .done(par_reset4_done)
  );
  
  std_reg #(1) par_done_reg15 (
      .in(par_done_reg15_in),
      .write_en(par_done_reg15_write_en),
      .clk(clk),
      .out(par_done_reg15_out),
      .done(par_done_reg15_done)
  );
  
  std_reg #(1) par_done_reg16 (
      .in(par_done_reg16_in),
      .write_en(par_done_reg16_write_en),
      .clk(clk),
      .out(par_done_reg16_out),
      .done(par_done_reg16_done)
  );
  
  std_reg #(1) par_done_reg17 (
      .in(par_done_reg17_in),
      .write_en(par_done_reg17_write_en),
      .clk(clk),
      .out(par_done_reg17_out),
      .done(par_done_reg17_done)
  );
  
  std_reg #(1) par_done_reg18 (
      .in(par_done_reg18_in),
      .write_en(par_done_reg18_write_en),
      .clk(clk),
      .out(par_done_reg18_out),
      .done(par_done_reg18_done)
  );
  
  std_reg #(1) par_done_reg19 (
      .in(par_done_reg19_in),
      .write_en(par_done_reg19_write_en),
      .clk(clk),
      .out(par_done_reg19_out),
      .done(par_done_reg19_done)
  );
  
  std_reg #(1) par_done_reg20 (
      .in(par_done_reg20_in),
      .write_en(par_done_reg20_write_en),
      .clk(clk),
      .out(par_done_reg20_out),
      .done(par_done_reg20_done)
  );
  
  std_reg #(1) par_reset5 (
      .in(par_reset5_in),
      .write_en(par_reset5_write_en),
      .clk(clk),
      .out(par_reset5_out),
      .done(par_reset5_done)
  );
  
  std_reg #(1) par_done_reg21 (
      .in(par_done_reg21_in),
      .write_en(par_done_reg21_write_en),
      .clk(clk),
      .out(par_done_reg21_out),
      .done(par_done_reg21_done)
  );
  
  std_reg #(1) par_done_reg22 (
      .in(par_done_reg22_in),
      .write_en(par_done_reg22_write_en),
      .clk(clk),
      .out(par_done_reg22_out),
      .done(par_done_reg22_done)
  );
  
  std_reg #(1) par_done_reg23 (
      .in(par_done_reg23_in),
      .write_en(par_done_reg23_write_en),
      .clk(clk),
      .out(par_done_reg23_out),
      .done(par_done_reg23_done)
  );
  
  std_reg #(1) par_done_reg24 (
      .in(par_done_reg24_in),
      .write_en(par_done_reg24_write_en),
      .clk(clk),
      .out(par_done_reg24_out),
      .done(par_done_reg24_done)
  );
  
  std_reg #(1) par_done_reg25 (
      .in(par_done_reg25_in),
      .write_en(par_done_reg25_write_en),
      .clk(clk),
      .out(par_done_reg25_out),
      .done(par_done_reg25_done)
  );
  
  std_reg #(1) par_done_reg26 (
      .in(par_done_reg26_in),
      .write_en(par_done_reg26_write_en),
      .clk(clk),
      .out(par_done_reg26_out),
      .done(par_done_reg26_done)
  );
  
  std_reg #(1) par_done_reg27 (
      .in(par_done_reg27_in),
      .write_en(par_done_reg27_write_en),
      .clk(clk),
      .out(par_done_reg27_out),
      .done(par_done_reg27_done)
  );
  
  std_reg #(1) par_done_reg28 (
      .in(par_done_reg28_in),
      .write_en(par_done_reg28_write_en),
      .clk(clk),
      .out(par_done_reg28_out),
      .done(par_done_reg28_done)
  );
  
  std_reg #(1) par_done_reg29 (
      .in(par_done_reg29_in),
      .write_en(par_done_reg29_write_en),
      .clk(clk),
      .out(par_done_reg29_out),
      .done(par_done_reg29_done)
  );
  
  std_reg #(1) par_reset6 (
      .in(par_reset6_in),
      .write_en(par_reset6_write_en),
      .clk(clk),
      .out(par_reset6_out),
      .done(par_reset6_done)
  );
  
  std_reg #(1) par_done_reg30 (
      .in(par_done_reg30_in),
      .write_en(par_done_reg30_write_en),
      .clk(clk),
      .out(par_done_reg30_out),
      .done(par_done_reg30_done)
  );
  
  std_reg #(1) par_done_reg31 (
      .in(par_done_reg31_in),
      .write_en(par_done_reg31_write_en),
      .clk(clk),
      .out(par_done_reg31_out),
      .done(par_done_reg31_done)
  );
  
  std_reg #(1) par_done_reg32 (
      .in(par_done_reg32_in),
      .write_en(par_done_reg32_write_en),
      .clk(clk),
      .out(par_done_reg32_out),
      .done(par_done_reg32_done)
  );
  
  std_reg #(1) par_done_reg33 (
      .in(par_done_reg33_in),
      .write_en(par_done_reg33_write_en),
      .clk(clk),
      .out(par_done_reg33_out),
      .done(par_done_reg33_done)
  );
  
  std_reg #(1) par_done_reg34 (
      .in(par_done_reg34_in),
      .write_en(par_done_reg34_write_en),
      .clk(clk),
      .out(par_done_reg34_out),
      .done(par_done_reg34_done)
  );
  
  std_reg #(1) par_done_reg35 (
      .in(par_done_reg35_in),
      .write_en(par_done_reg35_write_en),
      .clk(clk),
      .out(par_done_reg35_out),
      .done(par_done_reg35_done)
  );
  
  std_reg #(1) par_done_reg36 (
      .in(par_done_reg36_in),
      .write_en(par_done_reg36_write_en),
      .clk(clk),
      .out(par_done_reg36_out),
      .done(par_done_reg36_done)
  );
  
  std_reg #(1) par_done_reg37 (
      .in(par_done_reg37_in),
      .write_en(par_done_reg37_write_en),
      .clk(clk),
      .out(par_done_reg37_out),
      .done(par_done_reg37_done)
  );
  
  std_reg #(1) par_done_reg38 (
      .in(par_done_reg38_in),
      .write_en(par_done_reg38_write_en),
      .clk(clk),
      .out(par_done_reg38_out),
      .done(par_done_reg38_done)
  );
  
  std_reg #(1) par_done_reg39 (
      .in(par_done_reg39_in),
      .write_en(par_done_reg39_write_en),
      .clk(clk),
      .out(par_done_reg39_out),
      .done(par_done_reg39_done)
  );
  
  std_reg #(1) par_done_reg40 (
      .in(par_done_reg40_in),
      .write_en(par_done_reg40_write_en),
      .clk(clk),
      .out(par_done_reg40_out),
      .done(par_done_reg40_done)
  );
  
  std_reg #(1) par_done_reg41 (
      .in(par_done_reg41_in),
      .write_en(par_done_reg41_write_en),
      .clk(clk),
      .out(par_done_reg41_out),
      .done(par_done_reg41_done)
  );
  
  std_reg #(1) par_reset7 (
      .in(par_reset7_in),
      .write_en(par_reset7_write_en),
      .clk(clk),
      .out(par_reset7_out),
      .done(par_reset7_done)
  );
  
  std_reg #(1) par_done_reg42 (
      .in(par_done_reg42_in),
      .write_en(par_done_reg42_write_en),
      .clk(clk),
      .out(par_done_reg42_out),
      .done(par_done_reg42_done)
  );
  
  std_reg #(1) par_done_reg43 (
      .in(par_done_reg43_in),
      .write_en(par_done_reg43_write_en),
      .clk(clk),
      .out(par_done_reg43_out),
      .done(par_done_reg43_done)
  );
  
  std_reg #(1) par_done_reg44 (
      .in(par_done_reg44_in),
      .write_en(par_done_reg44_write_en),
      .clk(clk),
      .out(par_done_reg44_out),
      .done(par_done_reg44_done)
  );
  
  std_reg #(1) par_done_reg45 (
      .in(par_done_reg45_in),
      .write_en(par_done_reg45_write_en),
      .clk(clk),
      .out(par_done_reg45_out),
      .done(par_done_reg45_done)
  );
  
  std_reg #(1) par_done_reg46 (
      .in(par_done_reg46_in),
      .write_en(par_done_reg46_write_en),
      .clk(clk),
      .out(par_done_reg46_out),
      .done(par_done_reg46_done)
  );
  
  std_reg #(1) par_done_reg47 (
      .in(par_done_reg47_in),
      .write_en(par_done_reg47_write_en),
      .clk(clk),
      .out(par_done_reg47_out),
      .done(par_done_reg47_done)
  );
  
  std_reg #(1) par_done_reg48 (
      .in(par_done_reg48_in),
      .write_en(par_done_reg48_write_en),
      .clk(clk),
      .out(par_done_reg48_out),
      .done(par_done_reg48_done)
  );
  
  std_reg #(1) par_done_reg49 (
      .in(par_done_reg49_in),
      .write_en(par_done_reg49_write_en),
      .clk(clk),
      .out(par_done_reg49_out),
      .done(par_done_reg49_done)
  );
  
  std_reg #(1) par_done_reg50 (
      .in(par_done_reg50_in),
      .write_en(par_done_reg50_write_en),
      .clk(clk),
      .out(par_done_reg50_out),
      .done(par_done_reg50_done)
  );
  
  std_reg #(1) par_done_reg51 (
      .in(par_done_reg51_in),
      .write_en(par_done_reg51_write_en),
      .clk(clk),
      .out(par_done_reg51_out),
      .done(par_done_reg51_done)
  );
  
  std_reg #(1) par_reset8 (
      .in(par_reset8_in),
      .write_en(par_reset8_write_en),
      .clk(clk),
      .out(par_reset8_out),
      .done(par_reset8_done)
  );
  
  std_reg #(1) par_done_reg52 (
      .in(par_done_reg52_in),
      .write_en(par_done_reg52_write_en),
      .clk(clk),
      .out(par_done_reg52_out),
      .done(par_done_reg52_done)
  );
  
  std_reg #(1) par_done_reg53 (
      .in(par_done_reg53_in),
      .write_en(par_done_reg53_write_en),
      .clk(clk),
      .out(par_done_reg53_out),
      .done(par_done_reg53_done)
  );
  
  std_reg #(1) par_done_reg54 (
      .in(par_done_reg54_in),
      .write_en(par_done_reg54_write_en),
      .clk(clk),
      .out(par_done_reg54_out),
      .done(par_done_reg54_done)
  );
  
  std_reg #(1) par_done_reg55 (
      .in(par_done_reg55_in),
      .write_en(par_done_reg55_write_en),
      .clk(clk),
      .out(par_done_reg55_out),
      .done(par_done_reg55_done)
  );
  
  std_reg #(1) par_done_reg56 (
      .in(par_done_reg56_in),
      .write_en(par_done_reg56_write_en),
      .clk(clk),
      .out(par_done_reg56_out),
      .done(par_done_reg56_done)
  );
  
  std_reg #(1) par_done_reg57 (
      .in(par_done_reg57_in),
      .write_en(par_done_reg57_write_en),
      .clk(clk),
      .out(par_done_reg57_out),
      .done(par_done_reg57_done)
  );
  
  std_reg #(1) par_done_reg58 (
      .in(par_done_reg58_in),
      .write_en(par_done_reg58_write_en),
      .clk(clk),
      .out(par_done_reg58_out),
      .done(par_done_reg58_done)
  );
  
  std_reg #(1) par_done_reg59 (
      .in(par_done_reg59_in),
      .write_en(par_done_reg59_write_en),
      .clk(clk),
      .out(par_done_reg59_out),
      .done(par_done_reg59_done)
  );
  
  std_reg #(1) par_done_reg60 (
      .in(par_done_reg60_in),
      .write_en(par_done_reg60_write_en),
      .clk(clk),
      .out(par_done_reg60_out),
      .done(par_done_reg60_done)
  );
  
  std_reg #(1) par_done_reg61 (
      .in(par_done_reg61_in),
      .write_en(par_done_reg61_write_en),
      .clk(clk),
      .out(par_done_reg61_out),
      .done(par_done_reg61_done)
  );
  
  std_reg #(1) par_done_reg62 (
      .in(par_done_reg62_in),
      .write_en(par_done_reg62_write_en),
      .clk(clk),
      .out(par_done_reg62_out),
      .done(par_done_reg62_done)
  );
  
  std_reg #(1) par_done_reg63 (
      .in(par_done_reg63_in),
      .write_en(par_done_reg63_write_en),
      .clk(clk),
      .out(par_done_reg63_out),
      .done(par_done_reg63_done)
  );
  
  std_reg #(1) par_done_reg64 (
      .in(par_done_reg64_in),
      .write_en(par_done_reg64_write_en),
      .clk(clk),
      .out(par_done_reg64_out),
      .done(par_done_reg64_done)
  );
  
  std_reg #(1) par_done_reg65 (
      .in(par_done_reg65_in),
      .write_en(par_done_reg65_write_en),
      .clk(clk),
      .out(par_done_reg65_out),
      .done(par_done_reg65_done)
  );
  
  std_reg #(1) par_reset9 (
      .in(par_reset9_in),
      .write_en(par_reset9_write_en),
      .clk(clk),
      .out(par_reset9_out),
      .done(par_reset9_done)
  );
  
  std_reg #(1) par_done_reg66 (
      .in(par_done_reg66_in),
      .write_en(par_done_reg66_write_en),
      .clk(clk),
      .out(par_done_reg66_out),
      .done(par_done_reg66_done)
  );
  
  std_reg #(1) par_done_reg67 (
      .in(par_done_reg67_in),
      .write_en(par_done_reg67_write_en),
      .clk(clk),
      .out(par_done_reg67_out),
      .done(par_done_reg67_done)
  );
  
  std_reg #(1) par_done_reg68 (
      .in(par_done_reg68_in),
      .write_en(par_done_reg68_write_en),
      .clk(clk),
      .out(par_done_reg68_out),
      .done(par_done_reg68_done)
  );
  
  std_reg #(1) par_done_reg69 (
      .in(par_done_reg69_in),
      .write_en(par_done_reg69_write_en),
      .clk(clk),
      .out(par_done_reg69_out),
      .done(par_done_reg69_done)
  );
  
  std_reg #(1) par_done_reg70 (
      .in(par_done_reg70_in),
      .write_en(par_done_reg70_write_en),
      .clk(clk),
      .out(par_done_reg70_out),
      .done(par_done_reg70_done)
  );
  
  std_reg #(1) par_done_reg71 (
      .in(par_done_reg71_in),
      .write_en(par_done_reg71_write_en),
      .clk(clk),
      .out(par_done_reg71_out),
      .done(par_done_reg71_done)
  );
  
  std_reg #(1) par_done_reg72 (
      .in(par_done_reg72_in),
      .write_en(par_done_reg72_write_en),
      .clk(clk),
      .out(par_done_reg72_out),
      .done(par_done_reg72_done)
  );
  
  std_reg #(1) par_done_reg73 (
      .in(par_done_reg73_in),
      .write_en(par_done_reg73_write_en),
      .clk(clk),
      .out(par_done_reg73_out),
      .done(par_done_reg73_done)
  );
  
  std_reg #(1) par_done_reg74 (
      .in(par_done_reg74_in),
      .write_en(par_done_reg74_write_en),
      .clk(clk),
      .out(par_done_reg74_out),
      .done(par_done_reg74_done)
  );
  
  std_reg #(1) par_reset10 (
      .in(par_reset10_in),
      .write_en(par_reset10_write_en),
      .clk(clk),
      .out(par_reset10_out),
      .done(par_reset10_done)
  );
  
  std_reg #(1) par_done_reg75 (
      .in(par_done_reg75_in),
      .write_en(par_done_reg75_write_en),
      .clk(clk),
      .out(par_done_reg75_out),
      .done(par_done_reg75_done)
  );
  
  std_reg #(1) par_done_reg76 (
      .in(par_done_reg76_in),
      .write_en(par_done_reg76_write_en),
      .clk(clk),
      .out(par_done_reg76_out),
      .done(par_done_reg76_done)
  );
  
  std_reg #(1) par_done_reg77 (
      .in(par_done_reg77_in),
      .write_en(par_done_reg77_write_en),
      .clk(clk),
      .out(par_done_reg77_out),
      .done(par_done_reg77_done)
  );
  
  std_reg #(1) par_done_reg78 (
      .in(par_done_reg78_in),
      .write_en(par_done_reg78_write_en),
      .clk(clk),
      .out(par_done_reg78_out),
      .done(par_done_reg78_done)
  );
  
  std_reg #(1) par_done_reg79 (
      .in(par_done_reg79_in),
      .write_en(par_done_reg79_write_en),
      .clk(clk),
      .out(par_done_reg79_out),
      .done(par_done_reg79_done)
  );
  
  std_reg #(1) par_done_reg80 (
      .in(par_done_reg80_in),
      .write_en(par_done_reg80_write_en),
      .clk(clk),
      .out(par_done_reg80_out),
      .done(par_done_reg80_done)
  );
  
  std_reg #(1) par_done_reg81 (
      .in(par_done_reg81_in),
      .write_en(par_done_reg81_write_en),
      .clk(clk),
      .out(par_done_reg81_out),
      .done(par_done_reg81_done)
  );
  
  std_reg #(1) par_done_reg82 (
      .in(par_done_reg82_in),
      .write_en(par_done_reg82_write_en),
      .clk(clk),
      .out(par_done_reg82_out),
      .done(par_done_reg82_done)
  );
  
  std_reg #(1) par_done_reg83 (
      .in(par_done_reg83_in),
      .write_en(par_done_reg83_write_en),
      .clk(clk),
      .out(par_done_reg83_out),
      .done(par_done_reg83_done)
  );
  
  std_reg #(1) par_done_reg84 (
      .in(par_done_reg84_in),
      .write_en(par_done_reg84_write_en),
      .clk(clk),
      .out(par_done_reg84_out),
      .done(par_done_reg84_done)
  );
  
  std_reg #(1) par_done_reg85 (
      .in(par_done_reg85_in),
      .write_en(par_done_reg85_write_en),
      .clk(clk),
      .out(par_done_reg85_out),
      .done(par_done_reg85_done)
  );
  
  std_reg #(1) par_done_reg86 (
      .in(par_done_reg86_in),
      .write_en(par_done_reg86_write_en),
      .clk(clk),
      .out(par_done_reg86_out),
      .done(par_done_reg86_done)
  );
  
  std_reg #(1) par_reset11 (
      .in(par_reset11_in),
      .write_en(par_reset11_write_en),
      .clk(clk),
      .out(par_reset11_out),
      .done(par_reset11_done)
  );
  
  std_reg #(1) par_done_reg87 (
      .in(par_done_reg87_in),
      .write_en(par_done_reg87_write_en),
      .clk(clk),
      .out(par_done_reg87_out),
      .done(par_done_reg87_done)
  );
  
  std_reg #(1) par_done_reg88 (
      .in(par_done_reg88_in),
      .write_en(par_done_reg88_write_en),
      .clk(clk),
      .out(par_done_reg88_out),
      .done(par_done_reg88_done)
  );
  
  std_reg #(1) par_done_reg89 (
      .in(par_done_reg89_in),
      .write_en(par_done_reg89_write_en),
      .clk(clk),
      .out(par_done_reg89_out),
      .done(par_done_reg89_done)
  );
  
  std_reg #(1) par_done_reg90 (
      .in(par_done_reg90_in),
      .write_en(par_done_reg90_write_en),
      .clk(clk),
      .out(par_done_reg90_out),
      .done(par_done_reg90_done)
  );
  
  std_reg #(1) par_done_reg91 (
      .in(par_done_reg91_in),
      .write_en(par_done_reg91_write_en),
      .clk(clk),
      .out(par_done_reg91_out),
      .done(par_done_reg91_done)
  );
  
  std_reg #(1) par_done_reg92 (
      .in(par_done_reg92_in),
      .write_en(par_done_reg92_write_en),
      .clk(clk),
      .out(par_done_reg92_out),
      .done(par_done_reg92_done)
  );
  
  std_reg #(1) par_reset12 (
      .in(par_reset12_in),
      .write_en(par_reset12_write_en),
      .clk(clk),
      .out(par_reset12_out),
      .done(par_reset12_done)
  );
  
  std_reg #(1) par_done_reg93 (
      .in(par_done_reg93_in),
      .write_en(par_done_reg93_write_en),
      .clk(clk),
      .out(par_done_reg93_out),
      .done(par_done_reg93_done)
  );
  
  std_reg #(1) par_done_reg94 (
      .in(par_done_reg94_in),
      .write_en(par_done_reg94_write_en),
      .clk(clk),
      .out(par_done_reg94_out),
      .done(par_done_reg94_done)
  );
  
  std_reg #(1) par_done_reg95 (
      .in(par_done_reg95_in),
      .write_en(par_done_reg95_write_en),
      .clk(clk),
      .out(par_done_reg95_out),
      .done(par_done_reg95_done)
  );
  
  std_reg #(1) par_done_reg96 (
      .in(par_done_reg96_in),
      .write_en(par_done_reg96_write_en),
      .clk(clk),
      .out(par_done_reg96_out),
      .done(par_done_reg96_done)
  );
  
  std_reg #(1) par_done_reg97 (
      .in(par_done_reg97_in),
      .write_en(par_done_reg97_write_en),
      .clk(clk),
      .out(par_done_reg97_out),
      .done(par_done_reg97_done)
  );
  
  std_reg #(1) par_done_reg98 (
      .in(par_done_reg98_in),
      .write_en(par_done_reg98_write_en),
      .clk(clk),
      .out(par_done_reg98_out),
      .done(par_done_reg98_done)
  );
  
  std_reg #(1) par_reset13 (
      .in(par_reset13_in),
      .write_en(par_reset13_write_en),
      .clk(clk),
      .out(par_reset13_out),
      .done(par_reset13_done)
  );
  
  std_reg #(1) par_done_reg99 (
      .in(par_done_reg99_in),
      .write_en(par_done_reg99_write_en),
      .clk(clk),
      .out(par_done_reg99_out),
      .done(par_done_reg99_done)
  );
  
  std_reg #(1) par_done_reg100 (
      .in(par_done_reg100_in),
      .write_en(par_done_reg100_write_en),
      .clk(clk),
      .out(par_done_reg100_out),
      .done(par_done_reg100_done)
  );
  
  std_reg #(1) par_done_reg101 (
      .in(par_done_reg101_in),
      .write_en(par_done_reg101_write_en),
      .clk(clk),
      .out(par_done_reg101_out),
      .done(par_done_reg101_done)
  );
  
  std_reg #(1) par_reset14 (
      .in(par_reset14_in),
      .write_en(par_reset14_write_en),
      .clk(clk),
      .out(par_reset14_out),
      .done(par_reset14_done)
  );
  
  std_reg #(1) par_done_reg102 (
      .in(par_done_reg102_in),
      .write_en(par_done_reg102_write_en),
      .clk(clk),
      .out(par_done_reg102_out),
      .done(par_done_reg102_done)
  );
  
  std_reg #(1) par_done_reg103 (
      .in(par_done_reg103_in),
      .write_en(par_done_reg103_write_en),
      .clk(clk),
      .out(par_done_reg103_out),
      .done(par_done_reg103_done)
  );
  
  std_reg #(1) par_reset15 (
      .in(par_reset15_in),
      .write_en(par_reset15_write_en),
      .clk(clk),
      .out(par_reset15_out),
      .done(par_reset15_done)
  );
  
  std_reg #(1) par_done_reg104 (
      .in(par_done_reg104_in),
      .write_en(par_done_reg104_write_en),
      .clk(clk),
      .out(par_done_reg104_out),
      .done(par_done_reg104_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign done = (fsm0_out == 32'd25) ? 1'd1 : '0;
  assign out_mem_addr0 = (fsm0_out == 32'd22 & !out_mem_done & go | fsm0_out == 32'd23 & !out_mem_done & go | fsm0_out == 32'd24 & !out_mem_done & go) ? 2'd2 : (fsm0_out == 32'd16 & !out_mem_done & go | fsm0_out == 32'd17 & !out_mem_done & go | fsm0_out == 32'd18 & !out_mem_done & go) ? 2'd0 : (fsm0_out == 32'd19 & !out_mem_done & go | fsm0_out == 32'd20 & !out_mem_done & go | fsm0_out == 32'd21 & !out_mem_done & go) ? 2'd1 : '0;
  assign out_mem_addr1 = (fsm0_out == 32'd18 & !out_mem_done & go | fsm0_out == 32'd21 & !out_mem_done & go | fsm0_out == 32'd24 & !out_mem_done & go) ? 2'd2 : (fsm0_out == 32'd16 & !out_mem_done & go | fsm0_out == 32'd19 & !out_mem_done & go | fsm0_out == 32'd22 & !out_mem_done & go) ? 2'd0 : (fsm0_out == 32'd17 & !out_mem_done & go | fsm0_out == 32'd20 & !out_mem_done & go | fsm0_out == 32'd23 & !out_mem_done & go) ? 2'd1 : '0;
  assign out_mem_write_data = (fsm0_out == 32'd24 & !out_mem_done & go) ? pe_22_out : (fsm0_out == 32'd23 & !out_mem_done & go) ? pe_21_out : (fsm0_out == 32'd22 & !out_mem_done & go) ? pe_20_out : (fsm0_out == 32'd21 & !out_mem_done & go) ? pe_12_out : (fsm0_out == 32'd20 & !out_mem_done & go) ? pe_11_out : (fsm0_out == 32'd19 & !out_mem_done & go) ? pe_10_out : (fsm0_out == 32'd18 & !out_mem_done & go) ? pe_02_out : (fsm0_out == 32'd17 & !out_mem_done & go) ? pe_01_out : (fsm0_out == 32'd16 & !out_mem_done & go) ? pe_00_out : '0;
  assign out_mem_write_en = (fsm0_out == 32'd16 & !out_mem_done & go | fsm0_out == 32'd17 & !out_mem_done & go | fsm0_out == 32'd18 & !out_mem_done & go | fsm0_out == 32'd19 & !out_mem_done & go | fsm0_out == 32'd20 & !out_mem_done & go | fsm0_out == 32'd21 & !out_mem_done & go | fsm0_out == 32'd22 & !out_mem_done & go | fsm0_out == 32'd23 & !out_mem_done & go | fsm0_out == 32'd24 & !out_mem_done & go) ? 1'd1 : '0;
  assign left_22_read_in = (!(par_done_reg86_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg98_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg103_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_21_write_out : '0;
  assign left_22_read_write_en = (!(par_done_reg86_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg98_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg103_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_22_read_in = (!(par_done_reg80_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg95_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg102_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_12_write_out : '0;
  assign top_22_read_write_en = (!(par_done_reg80_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg95_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg102_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_22_top = (!(par_done_reg92_out | pe_22_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg101_out | pe_22_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg104_out | pe_22_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_22_read_out : '0;
  assign pe_22_left = (!(par_done_reg92_out | pe_22_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg101_out | pe_22_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg104_out | pe_22_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_22_read_out : '0;
  assign pe_22_go = (!pe_22_done & (!(par_done_reg92_out | pe_22_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg101_out | pe_22_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg104_out | pe_22_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_21_write_in = (pe_21_done & (!(par_done_reg74_out | right_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg91_out | right_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg100_out | right_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_21_right : '0;
  assign right_21_write_write_en = (pe_21_done & (!(par_done_reg74_out | right_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg91_out | right_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg100_out | right_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_21_read_in = (!(par_done_reg65_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg85_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg97_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? right_20_write_out : '0;
  assign left_21_read_write_en = (!(par_done_reg65_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg85_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg97_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_21_read_in = (!(par_done_reg58_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg79_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg94_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? down_11_write_out : '0;
  assign top_21_read_write_en = (!(par_done_reg58_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg79_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg94_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_21_top = (!(par_done_reg74_out | right_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg91_out | right_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg100_out | right_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_21_read_out : '0;
  assign pe_21_left = (!(par_done_reg74_out | right_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg91_out | right_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg100_out | right_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_21_read_out : '0;
  assign pe_21_go = (!pe_21_done & (!(par_done_reg74_out | right_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg91_out | right_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg100_out | right_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_20_write_in = (pe_20_done & (!(par_done_reg51_out | right_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg73_out | right_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg90_out | right_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_20_right : '0;
  assign right_20_write_write_en = (pe_20_done & (!(par_done_reg51_out | right_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg73_out | right_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg90_out | right_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign left_20_read_in = (!(par_done_reg41_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg84_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? l2_read_data : '0;
  assign left_20_read_write_en = (!(par_done_reg41_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg84_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign top_20_read_in = (!(par_done_reg35_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg57_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg78_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? down_10_write_out : '0;
  assign top_20_read_write_en = (!(par_done_reg35_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg57_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg78_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign pe_20_top = (!(par_done_reg51_out | right_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg73_out | right_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg90_out | right_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? top_20_read_out : '0;
  assign pe_20_left = (!(par_done_reg51_out | right_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg73_out | right_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg90_out | right_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? left_20_read_out : '0;
  assign pe_20_go = (!pe_20_done & (!(par_done_reg51_out | right_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg73_out | right_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg90_out | right_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign down_12_write_in = (pe_12_done & (!(par_done_reg72_out | down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg89_out | down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg99_out | down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_12_down : '0;
  assign down_12_write_write_en = (pe_12_done & (!(par_done_reg72_out | down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg89_out | down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg99_out | down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_12_read_in = (!(par_done_reg63_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg83_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg96_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? right_11_write_out : '0;
  assign left_12_read_write_en = (!(par_done_reg63_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg83_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg96_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_12_read_in = (!(par_done_reg56_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg77_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg93_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? down_02_write_out : '0;
  assign top_12_read_write_en = (!(par_done_reg56_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg77_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg93_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_12_top = (!(par_done_reg72_out | down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg89_out | down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg99_out | down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_12_read_out : '0;
  assign pe_12_left = (!(par_done_reg72_out | down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg89_out | down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg99_out | down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_12_read_out : '0;
  assign pe_12_go = (!pe_12_done & (!(par_done_reg72_out | down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg89_out | down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg99_out | down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign down_11_write_in = (pe_11_done & (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_11_down : '0;
  assign down_11_write_write_en = (pe_11_done & (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign right_11_write_in = (pe_11_done & (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_11_right : '0;
  assign right_11_write_write_en = (pe_11_done & (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign left_11_read_in = (!(par_done_reg40_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg82_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? right_10_write_out : '0;
  assign left_11_read_write_en = (!(par_done_reg40_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg82_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign top_11_read_in = (!(par_done_reg34_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg55_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg76_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? down_01_write_out : '0;
  assign top_11_read_write_en = (!(par_done_reg34_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg55_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg76_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign pe_11_top = (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? top_11_read_out : '0;
  assign pe_11_left = (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? left_11_read_out : '0;
  assign pe_11_go = (!pe_11_done & (!(par_done_reg50_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg71_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg88_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign down_10_write_in = (pe_10_done & (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? pe_10_down : '0;
  assign down_10_write_write_en = (pe_10_done & (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign right_10_write_in = (pe_10_done & (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? pe_10_right : '0;
  assign right_10_write_write_en = (pe_10_done & (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign left_10_read_in = (!(par_done_reg20_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg61_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? l1_read_data : '0;
  assign left_10_read_write_en = (!(par_done_reg20_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg61_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign top_10_read_in = (!(par_done_reg17_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg33_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg54_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? down_00_write_out : '0;
  assign top_10_read_write_en = (!(par_done_reg17_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg33_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg54_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign pe_10_top = (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? top_10_read_out : '0;
  assign pe_10_left = (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? left_10_read_out : '0;
  assign pe_10_go = (!pe_10_done & (!(par_done_reg29_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg70_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign down_02_write_in = (pe_02_done & (!(par_done_reg48_out | down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg69_out | down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg87_out | down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_02_down : '0;
  assign down_02_write_write_en = (pe_02_done & (!(par_done_reg48_out | down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg69_out | down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg87_out | down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign left_02_read_in = (!(par_done_reg38_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg81_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? right_01_write_out : '0;
  assign left_02_read_write_en = (!(par_done_reg38_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg81_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign top_02_read_in = (!(par_done_reg32_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg53_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg75_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? t2_read_data : '0;
  assign top_02_read_write_en = (!(par_done_reg32_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg53_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg75_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign pe_02_top = (!(par_done_reg48_out | down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg69_out | down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg87_out | down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? top_02_read_out : '0;
  assign pe_02_left = (!(par_done_reg48_out | down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg69_out | down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg87_out | down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? left_02_read_out : '0;
  assign pe_02_go = (!pe_02_done & (!(par_done_reg48_out | down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg69_out | down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg87_out | down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign down_01_write_in = (pe_01_done & (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? pe_01_down : '0;
  assign down_01_write_write_en = (pe_01_done & (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign right_01_write_in = (pe_01_done & (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? pe_01_right : '0;
  assign right_01_write_write_en = (pe_01_done & (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign left_01_read_in = (!(par_done_reg19_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg59_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? right_00_write_out : '0;
  assign left_01_read_write_en = (!(par_done_reg19_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg59_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign top_01_read_in = (!(par_done_reg16_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg31_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg52_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? t1_read_data : '0;
  assign top_01_read_write_en = (!(par_done_reg16_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg31_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg52_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign pe_01_top = (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? top_01_read_out : '0;
  assign pe_01_left = (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? left_01_read_out : '0;
  assign pe_01_go = (!pe_01_done & (!(par_done_reg28_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg68_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign down_00_write_in = (pe_00_done & (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go)) ? pe_00_down : '0;
  assign down_00_write_write_en = (pe_00_done & (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go)) ? 1'd1 : '0;
  assign right_00_write_in = (pe_00_done & (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go)) ? pe_00_right : '0;
  assign right_00_write_write_en = (pe_00_done & (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go)) ? 1'd1 : '0;
  assign left_00_read_in = (!(par_done_reg9_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg18_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg36_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go) ? l0_read_data : '0;
  assign left_00_read_write_en = (!(par_done_reg9_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg18_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg36_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign top_00_read_in = (!(par_done_reg8_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg15_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg30_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go) ? t0_read_data : '0;
  assign top_00_read_write_en = (!(par_done_reg8_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg15_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg30_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign pe_00_top = (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? top_00_read_out : '0;
  assign pe_00_left = (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? left_00_read_out : '0;
  assign pe_00_go = (!pe_00_done & (!(par_done_reg14_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go)) ? 1'd1 : '0;
  assign l2_addr0 = (!(par_done_reg41_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg84_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? l2_idx_out : '0;
  assign l2_add_left = (!(par_done_reg26_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg67_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 2'd1 : '0;
  assign l2_add_right = (!(par_done_reg26_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg67_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? l2_idx_out : '0;
  assign l2_idx_in = (!(par_done_reg26_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg67_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? l2_add_out : (!(par_done_reg5_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 2'd3 : '0;
  assign l2_idx_write_en = (!(par_done_reg5_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg26_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg67_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign l1_addr0 = (!(par_done_reg20_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg61_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? l1_idx_out : '0;
  assign l1_add_left = (!(par_done_reg13_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 2'd1 : '0;
  assign l1_add_right = (!(par_done_reg13_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? l1_idx_out : '0;
  assign l1_idx_in = (!(par_done_reg13_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? l1_add_out : (!(par_done_reg4_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 2'd3 : '0;
  assign l1_idx_write_en = (!(par_done_reg4_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg13_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign l0_addr0 = (!(par_done_reg9_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg18_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg36_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go) ? l0_idx_out : '0;
  assign l0_add_left = (!(par_done_reg7_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg22_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? 2'd1 : '0;
  assign l0_add_right = (!(par_done_reg7_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg22_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? l0_idx_out : '0;
  assign l0_idx_in = (!(par_done_reg7_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg22_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? l0_add_out : (!(par_done_reg3_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 2'd3 : '0;
  assign l0_idx_write_en = (!(par_done_reg3_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg7_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg11_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg22_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign t2_addr0 = (!(par_done_reg32_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg53_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg75_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? t2_idx_out : '0;
  assign t2_add_left = (!(par_done_reg24_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg43_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg66_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 2'd1 : '0;
  assign t2_add_right = (!(par_done_reg24_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg43_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg66_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? t2_idx_out : '0;
  assign t2_idx_in = (!(par_done_reg24_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg43_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg66_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? t2_add_out : (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 2'd3 : '0;
  assign t2_idx_write_en = (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg24_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg43_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg66_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign t1_addr0 = (!(par_done_reg16_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg31_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg52_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? t1_idx_out : '0;
  assign t1_add_left = (!(par_done_reg12_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg42_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 2'd1 : '0;
  assign t1_add_right = (!(par_done_reg12_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg42_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? t1_idx_out : '0;
  assign t1_idx_in = (!(par_done_reg12_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg42_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? t1_add_out : (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 2'd3 : '0;
  assign t1_idx_write_en = (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg12_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg42_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign t0_addr0 = (!(par_done_reg8_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg15_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg30_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go) ? t0_idx_out : '0;
  assign t0_add_left = (!(par_done_reg6_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg21_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? 2'd1 : '0;
  assign t0_add_right = (!(par_done_reg6_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg21_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? t0_idx_out : '0;
  assign t0_idx_in = (!(par_done_reg6_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg21_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? t0_add_out : (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 2'd3 : '0;
  assign t0_idx_write_en = (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg6_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg10_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg21_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_reset0_in = par_reset0_out ? 1'd0 : (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_reset0_write_en = (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg0_in = par_reset0_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg0_write_en = (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg1_in = par_reset0_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg1_write_en = (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg2_in = par_reset0_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg2_write_en = (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg3_in = par_reset0_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg3_write_en = (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg4_in = par_reset0_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg4_write_en = (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg5_in = par_reset0_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg5_write_en = (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_reset1_in = par_reset1_out ? 1'd0 : (par_done_reg6_out & par_done_reg7_out & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_reset1_write_en = (par_done_reg6_out & par_done_reg7_out & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg6_in = par_reset1_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg6_write_en = (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg7_in = par_reset1_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg7_write_en = (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_reset2_in = par_reset2_out ? 1'd0 : (par_done_reg8_out & par_done_reg9_out & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_reset2_write_en = (par_done_reg8_out & par_done_reg9_out & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg8_in = par_reset2_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg8_write_en = (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg9_in = par_reset2_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg9_write_en = (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_reset3_in = par_reset3_out ? 1'd0 : (par_done_reg10_out & par_done_reg11_out & par_done_reg12_out & par_done_reg13_out & par_done_reg14_out & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_reset3_write_en = (par_done_reg10_out & par_done_reg11_out & par_done_reg12_out & par_done_reg13_out & par_done_reg14_out & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg10_in = par_reset3_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg10_write_en = (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg11_in = par_reset3_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg11_write_en = (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg12_in = par_reset3_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg12_write_en = (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg13_in = par_reset3_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg13_write_en = (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg14_in = par_reset3_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg14_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_reset4_in = par_reset4_out ? 1'd0 : (par_done_reg15_out & par_done_reg16_out & par_done_reg17_out & par_done_reg18_out & par_done_reg19_out & par_done_reg20_out & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_reset4_write_en = (par_done_reg15_out & par_done_reg16_out & par_done_reg17_out & par_done_reg18_out & par_done_reg19_out & par_done_reg20_out & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg15_in = par_reset4_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg15_write_en = (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg16_in = par_reset4_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg16_write_en = (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg17_in = par_reset4_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg17_write_en = (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg18_in = par_reset4_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg18_write_en = (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg19_in = par_reset4_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg19_write_en = (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg20_in = par_reset4_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg20_write_en = (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_reset5_in = par_reset5_out ? 1'd0 : (par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_reset5_write_en = (par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg21_in = par_reset5_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg21_write_en = (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg22_in = par_reset5_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg22_write_en = (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg23_in = par_reset5_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg23_write_en = (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg24_in = par_reset5_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg24_write_en = (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg25_in = par_reset5_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg25_write_en = (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg26_in = par_reset5_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg26_write_en = (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg27_in = par_reset5_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg27_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg28_in = par_reset5_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg28_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg29_in = par_reset5_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg29_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_reset6_in = par_reset6_out ? 1'd0 : (par_done_reg30_out & par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_reset6_write_en = (par_done_reg30_out & par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg30_in = par_reset6_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg30_write_en = (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg31_in = par_reset6_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg31_write_en = (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg32_in = par_reset6_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg32_write_en = (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg33_in = par_reset6_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg33_write_en = (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg34_in = par_reset6_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg34_write_en = (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg35_in = par_reset6_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg35_write_en = (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg36_in = par_reset6_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg36_write_en = (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg37_in = par_reset6_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg37_write_en = (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg38_in = par_reset6_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg38_write_en = (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg39_in = par_reset6_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg39_write_en = (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg40_in = par_reset6_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg40_write_en = (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg41_in = par_reset6_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg41_write_en = (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_reset7_in = par_reset7_out ? 1'd0 : (par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_reset7_write_en = (par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg42_in = par_reset7_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg42_write_en = (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg43_in = par_reset7_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg43_write_en = (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg44_in = par_reset7_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg44_write_en = (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg45_in = par_reset7_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg45_write_en = (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg46_in = par_reset7_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg46_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg47_in = par_reset7_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg47_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg48_in = par_reset7_out ? 1'd0 : (down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg48_write_en = (down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg49_in = par_reset7_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg49_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg50_in = par_reset7_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg50_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg51_in = par_reset7_out ? 1'd0 : (right_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg51_write_en = (right_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_reset8_in = par_reset8_out ? 1'd0 : (par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_reset8_write_en = (par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg52_in = par_reset8_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg52_write_en = (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg53_in = par_reset8_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg53_write_en = (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg54_in = par_reset8_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg54_write_en = (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg55_in = par_reset8_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg55_write_en = (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg56_in = par_reset8_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg56_write_en = (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg57_in = par_reset8_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg57_write_en = (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg58_in = par_reset8_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg58_write_en = (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg59_in = par_reset8_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg59_write_en = (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg60_in = par_reset8_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg60_write_en = (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg61_in = par_reset8_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg61_write_en = (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg62_in = par_reset8_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg62_write_en = (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg63_in = par_reset8_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg63_write_en = (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg64_in = par_reset8_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg64_write_en = (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg65_in = par_reset8_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg65_write_en = (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_reset9_in = par_reset9_out ? 1'd0 : (par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_reset9_write_en = (par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg66_in = par_reset9_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg66_write_en = (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg67_in = par_reset9_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg67_write_en = (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg68_in = par_reset9_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg68_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg69_in = par_reset9_out ? 1'd0 : (down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg69_write_en = (down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg70_in = par_reset9_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg70_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg71_in = par_reset9_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg71_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg72_in = par_reset9_out ? 1'd0 : (down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg72_write_en = (down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg73_in = par_reset9_out ? 1'd0 : (right_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg73_write_en = (right_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg74_in = par_reset9_out ? 1'd0 : (right_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg74_write_en = (right_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_reset10_in = par_reset10_out ? 1'd0 : (par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_reset10_write_en = (par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg75_in = par_reset10_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg75_write_en = (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg76_in = par_reset10_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg76_write_en = (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg77_in = par_reset10_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg77_write_en = (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg78_in = par_reset10_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg78_write_en = (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg79_in = par_reset10_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg79_write_en = (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg80_in = par_reset10_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg80_write_en = (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg81_in = par_reset10_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg81_write_en = (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg82_in = par_reset10_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg82_write_en = (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg83_in = par_reset10_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg83_write_en = (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg84_in = par_reset10_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg84_write_en = (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg85_in = par_reset10_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg85_write_en = (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg86_in = par_reset10_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg86_write_en = (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_reset11_in = par_reset11_out ? 1'd0 : (par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_reset11_write_en = (par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg87_in = par_reset11_out ? 1'd0 : (down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg87_write_en = (down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg88_in = par_reset11_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg88_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg89_in = par_reset11_out ? 1'd0 : (down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg89_write_en = (down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg90_in = par_reset11_out ? 1'd0 : (right_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg90_write_en = (right_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg91_in = par_reset11_out ? 1'd0 : (right_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg91_write_en = (right_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg92_in = par_reset11_out ? 1'd0 : (pe_22_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg92_write_en = (pe_22_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_reset12_in = par_reset12_out ? 1'd0 : (par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_reset12_write_en = (par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg93_in = par_reset12_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg93_write_en = (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg94_in = par_reset12_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg94_write_en = (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg95_in = par_reset12_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg95_write_en = (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg96_in = par_reset12_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg96_write_en = (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg97_in = par_reset12_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg97_write_en = (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg98_in = par_reset12_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg98_write_en = (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_reset13_in = par_reset13_out ? 1'd0 : (par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_reset13_write_en = (par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg99_in = par_reset13_out ? 1'd0 : (down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg99_write_en = (down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg100_in = par_reset13_out ? 1'd0 : (right_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg100_write_en = (right_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg101_in = par_reset13_out ? 1'd0 : (pe_22_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg101_write_en = (pe_22_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_reset14_in = par_reset14_out ? 1'd0 : (par_done_reg102_out & par_done_reg103_out & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_reset14_write_en = (par_done_reg102_out & par_done_reg103_out & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg102_in = par_reset14_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg102_write_en = (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg103_in = par_reset14_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg103_write_en = (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_reset15_in = par_reset15_out ? 1'd0 : (par_done_reg104_out & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_reset15_write_en = (par_done_reg104_out & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg104_in = par_reset15_out ? 1'd0 : (pe_22_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg104_write_en = (pe_22_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd2 & par_reset2_out & go) ? 32'd3 : (fsm0_out == 32'd1 & par_reset1_out & go) ? 32'd2 : (fsm0_out == 32'd0 & par_reset0_out & go) ? 32'd1 : (fsm0_out == 32'd25) ? 32'd0 : (fsm0_out == 32'd24 & out_mem_done & go) ? 32'd25 : (fsm0_out == 32'd23 & out_mem_done & go) ? 32'd24 : (fsm0_out == 32'd22 & out_mem_done & go) ? 32'd23 : (fsm0_out == 32'd21 & out_mem_done & go) ? 32'd22 : (fsm0_out == 32'd20 & out_mem_done & go) ? 32'd21 : (fsm0_out == 32'd19 & out_mem_done & go) ? 32'd20 : (fsm0_out == 32'd18 & out_mem_done & go) ? 32'd19 : (fsm0_out == 32'd17 & out_mem_done & go) ? 32'd18 : (fsm0_out == 32'd16 & out_mem_done & go) ? 32'd17 : (fsm0_out == 32'd15 & par_reset15_out & go) ? 32'd16 : (fsm0_out == 32'd14 & par_reset14_out & go) ? 32'd15 : (fsm0_out == 32'd13 & par_reset13_out & go) ? 32'd14 : (fsm0_out == 32'd12 & par_reset12_out & go) ? 32'd13 : (fsm0_out == 32'd11 & par_reset11_out & go) ? 32'd12 : (fsm0_out == 32'd10 & par_reset10_out & go) ? 32'd11 : (fsm0_out == 32'd9 & par_reset9_out & go) ? 32'd10 : (fsm0_out == 32'd8 & par_reset8_out & go) ? 32'd9 : (fsm0_out == 32'd7 & par_reset7_out & go) ? 32'd8 : (fsm0_out == 32'd6 & par_reset6_out & go) ? 32'd7 : (fsm0_out == 32'd5 & par_reset5_out & go) ? 32'd6 : (fsm0_out == 32'd4 & par_reset4_out & go) ? 32'd5 : (fsm0_out == 32'd3 & par_reset3_out & go) ? 32'd4 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & par_reset0_out & go | fsm0_out == 32'd1 & par_reset1_out & go | fsm0_out == 32'd2 & par_reset2_out & go | fsm0_out == 32'd3 & par_reset3_out & go | fsm0_out == 32'd4 & par_reset4_out & go | fsm0_out == 32'd5 & par_reset5_out & go | fsm0_out == 32'd6 & par_reset6_out & go | fsm0_out == 32'd7 & par_reset7_out & go | fsm0_out == 32'd8 & par_reset8_out & go | fsm0_out == 32'd9 & par_reset9_out & go | fsm0_out == 32'd10 & par_reset10_out & go | fsm0_out == 32'd11 & par_reset11_out & go | fsm0_out == 32'd12 & par_reset12_out & go | fsm0_out == 32'd13 & par_reset13_out & go | fsm0_out == 32'd14 & par_reset14_out & go | fsm0_out == 32'd15 & par_reset15_out & go | fsm0_out == 32'd16 & out_mem_done & go | fsm0_out == 32'd17 & out_mem_done & go | fsm0_out == 32'd18 & out_mem_done & go | fsm0_out == 32'd19 & out_mem_done & go | fsm0_out == 32'd20 & out_mem_done & go | fsm0_out == 32'd21 & out_mem_done & go | fsm0_out == 32'd22 & out_mem_done & go | fsm0_out == 32'd23 & out_mem_done & go | fsm0_out == 32'd24 & out_mem_done & go | fsm0_out == 32'd25) ? 1'd1 : '0;
endmodule // end main