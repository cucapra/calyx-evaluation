/* verilator lint_off WIDTH */
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule

module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule

module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

// Component Signature
module mac_pe (
      input wire [31:0] top,
      input wire [31:0] left,
      input wire go,
      input wire clk,
      output wire [31:0] down,
      output wire [31:0] right,
      output wire [31:0] out,
      output wire done
  );
  
  // Structure wire declarations
  wire [31:0] mul_left;
  wire [31:0] mul_right;
  wire mul_go;
  wire mul_clk;
  wire [31:0] mul_out;
  wire mul_done;
  wire [31:0] add_left;
  wire [31:0] add_right;
  wire [31:0] add_out;
  wire [31:0] mul_reg_in;
  wire mul_reg_write_en;
  wire mul_reg_clk;
  wire [31:0] mul_reg_out;
  wire mul_reg_done;
  wire [31:0] acc_in;
  wire acc_write_en;
  wire acc_clk;
  wire [31:0] acc_out;
  wire acc_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_mult_pipe #(32) mul (
      .left(mul_left),
      .right(mul_right),
      .go(mul_go),
      .clk(clk),
      .out(mul_out),
      .done(mul_done)
  );
  
  std_add #(32) add (
      .left(add_left),
      .right(add_right),
      .out(add_out)
  );
  
  std_reg #(32) mul_reg (
      .in(mul_reg_in),
      .write_en(mul_reg_write_en),
      .clk(clk),
      .out(mul_reg_out),
      .done(mul_reg_done)
  );
  
  std_reg #(32) acc (
      .in(acc_in),
      .write_en(acc_write_en),
      .clk(clk),
      .out(acc_out),
      .done(acc_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign down = top;
  assign right = left;
  assign out = acc_out;
  assign done = (fsm0_out == 32'd2) ? 1'd1 : '0;
  assign mul_left = (fsm0_out == 32'd0 & !mul_reg_done & go) ? top : '0;
  assign mul_right = (fsm0_out == 32'd0 & !mul_reg_done & go) ? left : '0;
  assign mul_go = (!mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign add_left = (fsm0_out == 32'd1 & !acc_done & go) ? acc_out : '0;
  assign add_right = (fsm0_out == 32'd1 & !acc_done & go) ? mul_reg_out : '0;
  assign mul_reg_in = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? mul_out : '0;
  assign mul_reg_write_en = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign acc_in = (fsm0_out == 32'd1 & !acc_done & go) ? add_out : '0;
  assign acc_write_en = (fsm0_out == 32'd1 & !acc_done & go) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd1 & acc_done & go) ? 32'd2 : (fsm0_out == 32'd0 & mul_reg_done & go) ? 32'd1 : (fsm0_out == 32'd2) ? 32'd0 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & mul_reg_done & go | fsm0_out == 32'd1 & acc_done & go | fsm0_out == 32'd2) ? 1'd1 : '0;
endmodule // end mac_pe
// Component Signature
module main (
      input wire go,
      input wire clk,
      input wire [31:0] out_mem_read_data,
      input wire out_mem_done,
      output wire done,
      output wire [2:0] out_mem_addr0,
      output wire [2:0] out_mem_addr1,
      output wire [31:0] out_mem_write_data,
      output wire out_mem_write_en
  );
  
  // Structure wire declarations
  wire [31:0] left_33_read_in;
  wire left_33_read_write_en;
  wire left_33_read_clk;
  wire [31:0] left_33_read_out;
  wire left_33_read_done;
  wire [31:0] top_33_read_in;
  wire top_33_read_write_en;
  wire top_33_read_clk;
  wire [31:0] top_33_read_out;
  wire top_33_read_done;
  wire [31:0] pe_33_top;
  wire [31:0] pe_33_left;
  wire pe_33_go;
  wire pe_33_clk;
  wire [31:0] pe_33_down;
  wire [31:0] pe_33_right;
  wire [31:0] pe_33_out;
  wire pe_33_done;
  wire [31:0] right_32_write_in;
  wire right_32_write_write_en;
  wire right_32_write_clk;
  wire [31:0] right_32_write_out;
  wire right_32_write_done;
  wire [31:0] left_32_read_in;
  wire left_32_read_write_en;
  wire left_32_read_clk;
  wire [31:0] left_32_read_out;
  wire left_32_read_done;
  wire [31:0] top_32_read_in;
  wire top_32_read_write_en;
  wire top_32_read_clk;
  wire [31:0] top_32_read_out;
  wire top_32_read_done;
  wire [31:0] pe_32_top;
  wire [31:0] pe_32_left;
  wire pe_32_go;
  wire pe_32_clk;
  wire [31:0] pe_32_down;
  wire [31:0] pe_32_right;
  wire [31:0] pe_32_out;
  wire pe_32_done;
  wire [31:0] right_31_write_in;
  wire right_31_write_write_en;
  wire right_31_write_clk;
  wire [31:0] right_31_write_out;
  wire right_31_write_done;
  wire [31:0] left_31_read_in;
  wire left_31_read_write_en;
  wire left_31_read_clk;
  wire [31:0] left_31_read_out;
  wire left_31_read_done;
  wire [31:0] top_31_read_in;
  wire top_31_read_write_en;
  wire top_31_read_clk;
  wire [31:0] top_31_read_out;
  wire top_31_read_done;
  wire [31:0] pe_31_top;
  wire [31:0] pe_31_left;
  wire pe_31_go;
  wire pe_31_clk;
  wire [31:0] pe_31_down;
  wire [31:0] pe_31_right;
  wire [31:0] pe_31_out;
  wire pe_31_done;
  wire [31:0] right_30_write_in;
  wire right_30_write_write_en;
  wire right_30_write_clk;
  wire [31:0] right_30_write_out;
  wire right_30_write_done;
  wire [31:0] left_30_read_in;
  wire left_30_read_write_en;
  wire left_30_read_clk;
  wire [31:0] left_30_read_out;
  wire left_30_read_done;
  wire [31:0] top_30_read_in;
  wire top_30_read_write_en;
  wire top_30_read_clk;
  wire [31:0] top_30_read_out;
  wire top_30_read_done;
  wire [31:0] pe_30_top;
  wire [31:0] pe_30_left;
  wire pe_30_go;
  wire pe_30_clk;
  wire [31:0] pe_30_down;
  wire [31:0] pe_30_right;
  wire [31:0] pe_30_out;
  wire pe_30_done;
  wire [31:0] down_23_write_in;
  wire down_23_write_write_en;
  wire down_23_write_clk;
  wire [31:0] down_23_write_out;
  wire down_23_write_done;
  wire [31:0] left_23_read_in;
  wire left_23_read_write_en;
  wire left_23_read_clk;
  wire [31:0] left_23_read_out;
  wire left_23_read_done;
  wire [31:0] top_23_read_in;
  wire top_23_read_write_en;
  wire top_23_read_clk;
  wire [31:0] top_23_read_out;
  wire top_23_read_done;
  wire [31:0] pe_23_top;
  wire [31:0] pe_23_left;
  wire pe_23_go;
  wire pe_23_clk;
  wire [31:0] pe_23_down;
  wire [31:0] pe_23_right;
  wire [31:0] pe_23_out;
  wire pe_23_done;
  wire [31:0] down_22_write_in;
  wire down_22_write_write_en;
  wire down_22_write_clk;
  wire [31:0] down_22_write_out;
  wire down_22_write_done;
  wire [31:0] right_22_write_in;
  wire right_22_write_write_en;
  wire right_22_write_clk;
  wire [31:0] right_22_write_out;
  wire right_22_write_done;
  wire [31:0] left_22_read_in;
  wire left_22_read_write_en;
  wire left_22_read_clk;
  wire [31:0] left_22_read_out;
  wire left_22_read_done;
  wire [31:0] top_22_read_in;
  wire top_22_read_write_en;
  wire top_22_read_clk;
  wire [31:0] top_22_read_out;
  wire top_22_read_done;
  wire [31:0] pe_22_top;
  wire [31:0] pe_22_left;
  wire pe_22_go;
  wire pe_22_clk;
  wire [31:0] pe_22_down;
  wire [31:0] pe_22_right;
  wire [31:0] pe_22_out;
  wire pe_22_done;
  wire [31:0] down_21_write_in;
  wire down_21_write_write_en;
  wire down_21_write_clk;
  wire [31:0] down_21_write_out;
  wire down_21_write_done;
  wire [31:0] right_21_write_in;
  wire right_21_write_write_en;
  wire right_21_write_clk;
  wire [31:0] right_21_write_out;
  wire right_21_write_done;
  wire [31:0] left_21_read_in;
  wire left_21_read_write_en;
  wire left_21_read_clk;
  wire [31:0] left_21_read_out;
  wire left_21_read_done;
  wire [31:0] top_21_read_in;
  wire top_21_read_write_en;
  wire top_21_read_clk;
  wire [31:0] top_21_read_out;
  wire top_21_read_done;
  wire [31:0] pe_21_top;
  wire [31:0] pe_21_left;
  wire pe_21_go;
  wire pe_21_clk;
  wire [31:0] pe_21_down;
  wire [31:0] pe_21_right;
  wire [31:0] pe_21_out;
  wire pe_21_done;
  wire [31:0] down_20_write_in;
  wire down_20_write_write_en;
  wire down_20_write_clk;
  wire [31:0] down_20_write_out;
  wire down_20_write_done;
  wire [31:0] right_20_write_in;
  wire right_20_write_write_en;
  wire right_20_write_clk;
  wire [31:0] right_20_write_out;
  wire right_20_write_done;
  wire [31:0] left_20_read_in;
  wire left_20_read_write_en;
  wire left_20_read_clk;
  wire [31:0] left_20_read_out;
  wire left_20_read_done;
  wire [31:0] top_20_read_in;
  wire top_20_read_write_en;
  wire top_20_read_clk;
  wire [31:0] top_20_read_out;
  wire top_20_read_done;
  wire [31:0] pe_20_top;
  wire [31:0] pe_20_left;
  wire pe_20_go;
  wire pe_20_clk;
  wire [31:0] pe_20_down;
  wire [31:0] pe_20_right;
  wire [31:0] pe_20_out;
  wire pe_20_done;
  wire [31:0] down_13_write_in;
  wire down_13_write_write_en;
  wire down_13_write_clk;
  wire [31:0] down_13_write_out;
  wire down_13_write_done;
  wire [31:0] left_13_read_in;
  wire left_13_read_write_en;
  wire left_13_read_clk;
  wire [31:0] left_13_read_out;
  wire left_13_read_done;
  wire [31:0] top_13_read_in;
  wire top_13_read_write_en;
  wire top_13_read_clk;
  wire [31:0] top_13_read_out;
  wire top_13_read_done;
  wire [31:0] pe_13_top;
  wire [31:0] pe_13_left;
  wire pe_13_go;
  wire pe_13_clk;
  wire [31:0] pe_13_down;
  wire [31:0] pe_13_right;
  wire [31:0] pe_13_out;
  wire pe_13_done;
  wire [31:0] down_12_write_in;
  wire down_12_write_write_en;
  wire down_12_write_clk;
  wire [31:0] down_12_write_out;
  wire down_12_write_done;
  wire [31:0] right_12_write_in;
  wire right_12_write_write_en;
  wire right_12_write_clk;
  wire [31:0] right_12_write_out;
  wire right_12_write_done;
  wire [31:0] left_12_read_in;
  wire left_12_read_write_en;
  wire left_12_read_clk;
  wire [31:0] left_12_read_out;
  wire left_12_read_done;
  wire [31:0] top_12_read_in;
  wire top_12_read_write_en;
  wire top_12_read_clk;
  wire [31:0] top_12_read_out;
  wire top_12_read_done;
  wire [31:0] pe_12_top;
  wire [31:0] pe_12_left;
  wire pe_12_go;
  wire pe_12_clk;
  wire [31:0] pe_12_down;
  wire [31:0] pe_12_right;
  wire [31:0] pe_12_out;
  wire pe_12_done;
  wire [31:0] down_11_write_in;
  wire down_11_write_write_en;
  wire down_11_write_clk;
  wire [31:0] down_11_write_out;
  wire down_11_write_done;
  wire [31:0] right_11_write_in;
  wire right_11_write_write_en;
  wire right_11_write_clk;
  wire [31:0] right_11_write_out;
  wire right_11_write_done;
  wire [31:0] left_11_read_in;
  wire left_11_read_write_en;
  wire left_11_read_clk;
  wire [31:0] left_11_read_out;
  wire left_11_read_done;
  wire [31:0] top_11_read_in;
  wire top_11_read_write_en;
  wire top_11_read_clk;
  wire [31:0] top_11_read_out;
  wire top_11_read_done;
  wire [31:0] pe_11_top;
  wire [31:0] pe_11_left;
  wire pe_11_go;
  wire pe_11_clk;
  wire [31:0] pe_11_down;
  wire [31:0] pe_11_right;
  wire [31:0] pe_11_out;
  wire pe_11_done;
  wire [31:0] down_10_write_in;
  wire down_10_write_write_en;
  wire down_10_write_clk;
  wire [31:0] down_10_write_out;
  wire down_10_write_done;
  wire [31:0] right_10_write_in;
  wire right_10_write_write_en;
  wire right_10_write_clk;
  wire [31:0] right_10_write_out;
  wire right_10_write_done;
  wire [31:0] left_10_read_in;
  wire left_10_read_write_en;
  wire left_10_read_clk;
  wire [31:0] left_10_read_out;
  wire left_10_read_done;
  wire [31:0] top_10_read_in;
  wire top_10_read_write_en;
  wire top_10_read_clk;
  wire [31:0] top_10_read_out;
  wire top_10_read_done;
  wire [31:0] pe_10_top;
  wire [31:0] pe_10_left;
  wire pe_10_go;
  wire pe_10_clk;
  wire [31:0] pe_10_down;
  wire [31:0] pe_10_right;
  wire [31:0] pe_10_out;
  wire pe_10_done;
  wire [31:0] down_03_write_in;
  wire down_03_write_write_en;
  wire down_03_write_clk;
  wire [31:0] down_03_write_out;
  wire down_03_write_done;
  wire [31:0] left_03_read_in;
  wire left_03_read_write_en;
  wire left_03_read_clk;
  wire [31:0] left_03_read_out;
  wire left_03_read_done;
  wire [31:0] top_03_read_in;
  wire top_03_read_write_en;
  wire top_03_read_clk;
  wire [31:0] top_03_read_out;
  wire top_03_read_done;
  wire [31:0] pe_03_top;
  wire [31:0] pe_03_left;
  wire pe_03_go;
  wire pe_03_clk;
  wire [31:0] pe_03_down;
  wire [31:0] pe_03_right;
  wire [31:0] pe_03_out;
  wire pe_03_done;
  wire [31:0] down_02_write_in;
  wire down_02_write_write_en;
  wire down_02_write_clk;
  wire [31:0] down_02_write_out;
  wire down_02_write_done;
  wire [31:0] right_02_write_in;
  wire right_02_write_write_en;
  wire right_02_write_clk;
  wire [31:0] right_02_write_out;
  wire right_02_write_done;
  wire [31:0] left_02_read_in;
  wire left_02_read_write_en;
  wire left_02_read_clk;
  wire [31:0] left_02_read_out;
  wire left_02_read_done;
  wire [31:0] top_02_read_in;
  wire top_02_read_write_en;
  wire top_02_read_clk;
  wire [31:0] top_02_read_out;
  wire top_02_read_done;
  wire [31:0] pe_02_top;
  wire [31:0] pe_02_left;
  wire pe_02_go;
  wire pe_02_clk;
  wire [31:0] pe_02_down;
  wire [31:0] pe_02_right;
  wire [31:0] pe_02_out;
  wire pe_02_done;
  wire [31:0] down_01_write_in;
  wire down_01_write_write_en;
  wire down_01_write_clk;
  wire [31:0] down_01_write_out;
  wire down_01_write_done;
  wire [31:0] right_01_write_in;
  wire right_01_write_write_en;
  wire right_01_write_clk;
  wire [31:0] right_01_write_out;
  wire right_01_write_done;
  wire [31:0] left_01_read_in;
  wire left_01_read_write_en;
  wire left_01_read_clk;
  wire [31:0] left_01_read_out;
  wire left_01_read_done;
  wire [31:0] top_01_read_in;
  wire top_01_read_write_en;
  wire top_01_read_clk;
  wire [31:0] top_01_read_out;
  wire top_01_read_done;
  wire [31:0] pe_01_top;
  wire [31:0] pe_01_left;
  wire pe_01_go;
  wire pe_01_clk;
  wire [31:0] pe_01_down;
  wire [31:0] pe_01_right;
  wire [31:0] pe_01_out;
  wire pe_01_done;
  wire [31:0] down_00_write_in;
  wire down_00_write_write_en;
  wire down_00_write_clk;
  wire [31:0] down_00_write_out;
  wire down_00_write_done;
  wire [31:0] right_00_write_in;
  wire right_00_write_write_en;
  wire right_00_write_clk;
  wire [31:0] right_00_write_out;
  wire right_00_write_done;
  wire [31:0] left_00_read_in;
  wire left_00_read_write_en;
  wire left_00_read_clk;
  wire [31:0] left_00_read_out;
  wire left_00_read_done;
  wire [31:0] top_00_read_in;
  wire top_00_read_write_en;
  wire top_00_read_clk;
  wire [31:0] top_00_read_out;
  wire top_00_read_done;
  wire [31:0] pe_00_top;
  wire [31:0] pe_00_left;
  wire pe_00_go;
  wire pe_00_clk;
  wire [31:0] pe_00_down;
  wire [31:0] pe_00_right;
  wire [31:0] pe_00_out;
  wire pe_00_done;
  wire [2:0] l3_addr0;
  wire [31:0] l3_write_data;
  wire l3_write_en;
  wire l3_clk;
  wire [31:0] l3_read_data;
  wire l3_done;
  wire [2:0] l3_add_left;
  wire [2:0] l3_add_right;
  wire [2:0] l3_add_out;
  wire [2:0] l3_idx_in;
  wire l3_idx_write_en;
  wire l3_idx_clk;
  wire [2:0] l3_idx_out;
  wire l3_idx_done;
  wire [2:0] l2_addr0;
  wire [31:0] l2_write_data;
  wire l2_write_en;
  wire l2_clk;
  wire [31:0] l2_read_data;
  wire l2_done;
  wire [2:0] l2_add_left;
  wire [2:0] l2_add_right;
  wire [2:0] l2_add_out;
  wire [2:0] l2_idx_in;
  wire l2_idx_write_en;
  wire l2_idx_clk;
  wire [2:0] l2_idx_out;
  wire l2_idx_done;
  wire [2:0] l1_addr0;
  wire [31:0] l1_write_data;
  wire l1_write_en;
  wire l1_clk;
  wire [31:0] l1_read_data;
  wire l1_done;
  wire [2:0] l1_add_left;
  wire [2:0] l1_add_right;
  wire [2:0] l1_add_out;
  wire [2:0] l1_idx_in;
  wire l1_idx_write_en;
  wire l1_idx_clk;
  wire [2:0] l1_idx_out;
  wire l1_idx_done;
  wire [2:0] l0_addr0;
  wire [31:0] l0_write_data;
  wire l0_write_en;
  wire l0_clk;
  wire [31:0] l0_read_data;
  wire l0_done;
  wire [2:0] l0_add_left;
  wire [2:0] l0_add_right;
  wire [2:0] l0_add_out;
  wire [2:0] l0_idx_in;
  wire l0_idx_write_en;
  wire l0_idx_clk;
  wire [2:0] l0_idx_out;
  wire l0_idx_done;
  wire [2:0] t3_addr0;
  wire [31:0] t3_write_data;
  wire t3_write_en;
  wire t3_clk;
  wire [31:0] t3_read_data;
  wire t3_done;
  wire [2:0] t3_add_left;
  wire [2:0] t3_add_right;
  wire [2:0] t3_add_out;
  wire [2:0] t3_idx_in;
  wire t3_idx_write_en;
  wire t3_idx_clk;
  wire [2:0] t3_idx_out;
  wire t3_idx_done;
  wire [2:0] t2_addr0;
  wire [31:0] t2_write_data;
  wire t2_write_en;
  wire t2_clk;
  wire [31:0] t2_read_data;
  wire t2_done;
  wire [2:0] t2_add_left;
  wire [2:0] t2_add_right;
  wire [2:0] t2_add_out;
  wire [2:0] t2_idx_in;
  wire t2_idx_write_en;
  wire t2_idx_clk;
  wire [2:0] t2_idx_out;
  wire t2_idx_done;
  wire [2:0] t1_addr0;
  wire [31:0] t1_write_data;
  wire t1_write_en;
  wire t1_clk;
  wire [31:0] t1_read_data;
  wire t1_done;
  wire [2:0] t1_add_left;
  wire [2:0] t1_add_right;
  wire [2:0] t1_add_out;
  wire [2:0] t1_idx_in;
  wire t1_idx_write_en;
  wire t1_idx_clk;
  wire [2:0] t1_idx_out;
  wire t1_idx_done;
  wire [2:0] t0_addr0;
  wire [31:0] t0_write_data;
  wire t0_write_en;
  wire t0_clk;
  wire [31:0] t0_read_data;
  wire t0_done;
  wire [2:0] t0_add_left;
  wire [2:0] t0_add_right;
  wire [2:0] t0_add_out;
  wire [2:0] t0_idx_in;
  wire t0_idx_write_en;
  wire t0_idx_clk;
  wire [2:0] t0_idx_out;
  wire t0_idx_done;
  wire par_reset0_in;
  wire par_reset0_write_en;
  wire par_reset0_clk;
  wire par_reset0_out;
  wire par_reset0_done;
  wire par_done_reg0_in;
  wire par_done_reg0_write_en;
  wire par_done_reg0_clk;
  wire par_done_reg0_out;
  wire par_done_reg0_done;
  wire par_done_reg1_in;
  wire par_done_reg1_write_en;
  wire par_done_reg1_clk;
  wire par_done_reg1_out;
  wire par_done_reg1_done;
  wire par_done_reg2_in;
  wire par_done_reg2_write_en;
  wire par_done_reg2_clk;
  wire par_done_reg2_out;
  wire par_done_reg2_done;
  wire par_done_reg3_in;
  wire par_done_reg3_write_en;
  wire par_done_reg3_clk;
  wire par_done_reg3_out;
  wire par_done_reg3_done;
  wire par_done_reg4_in;
  wire par_done_reg4_write_en;
  wire par_done_reg4_clk;
  wire par_done_reg4_out;
  wire par_done_reg4_done;
  wire par_done_reg5_in;
  wire par_done_reg5_write_en;
  wire par_done_reg5_clk;
  wire par_done_reg5_out;
  wire par_done_reg5_done;
  wire par_done_reg6_in;
  wire par_done_reg6_write_en;
  wire par_done_reg6_clk;
  wire par_done_reg6_out;
  wire par_done_reg6_done;
  wire par_done_reg7_in;
  wire par_done_reg7_write_en;
  wire par_done_reg7_clk;
  wire par_done_reg7_out;
  wire par_done_reg7_done;
  wire par_reset1_in;
  wire par_reset1_write_en;
  wire par_reset1_clk;
  wire par_reset1_out;
  wire par_reset1_done;
  wire par_done_reg8_in;
  wire par_done_reg8_write_en;
  wire par_done_reg8_clk;
  wire par_done_reg8_out;
  wire par_done_reg8_done;
  wire par_done_reg9_in;
  wire par_done_reg9_write_en;
  wire par_done_reg9_clk;
  wire par_done_reg9_out;
  wire par_done_reg9_done;
  wire par_reset2_in;
  wire par_reset2_write_en;
  wire par_reset2_clk;
  wire par_reset2_out;
  wire par_reset2_done;
  wire par_done_reg10_in;
  wire par_done_reg10_write_en;
  wire par_done_reg10_clk;
  wire par_done_reg10_out;
  wire par_done_reg10_done;
  wire par_done_reg11_in;
  wire par_done_reg11_write_en;
  wire par_done_reg11_clk;
  wire par_done_reg11_out;
  wire par_done_reg11_done;
  wire par_reset3_in;
  wire par_reset3_write_en;
  wire par_reset3_clk;
  wire par_reset3_out;
  wire par_reset3_done;
  wire par_done_reg12_in;
  wire par_done_reg12_write_en;
  wire par_done_reg12_clk;
  wire par_done_reg12_out;
  wire par_done_reg12_done;
  wire par_done_reg13_in;
  wire par_done_reg13_write_en;
  wire par_done_reg13_clk;
  wire par_done_reg13_out;
  wire par_done_reg13_done;
  wire par_done_reg14_in;
  wire par_done_reg14_write_en;
  wire par_done_reg14_clk;
  wire par_done_reg14_out;
  wire par_done_reg14_done;
  wire par_done_reg15_in;
  wire par_done_reg15_write_en;
  wire par_done_reg15_clk;
  wire par_done_reg15_out;
  wire par_done_reg15_done;
  wire par_done_reg16_in;
  wire par_done_reg16_write_en;
  wire par_done_reg16_clk;
  wire par_done_reg16_out;
  wire par_done_reg16_done;
  wire par_reset4_in;
  wire par_reset4_write_en;
  wire par_reset4_clk;
  wire par_reset4_out;
  wire par_reset4_done;
  wire par_done_reg17_in;
  wire par_done_reg17_write_en;
  wire par_done_reg17_clk;
  wire par_done_reg17_out;
  wire par_done_reg17_done;
  wire par_done_reg18_in;
  wire par_done_reg18_write_en;
  wire par_done_reg18_clk;
  wire par_done_reg18_out;
  wire par_done_reg18_done;
  wire par_done_reg19_in;
  wire par_done_reg19_write_en;
  wire par_done_reg19_clk;
  wire par_done_reg19_out;
  wire par_done_reg19_done;
  wire par_done_reg20_in;
  wire par_done_reg20_write_en;
  wire par_done_reg20_clk;
  wire par_done_reg20_out;
  wire par_done_reg20_done;
  wire par_done_reg21_in;
  wire par_done_reg21_write_en;
  wire par_done_reg21_clk;
  wire par_done_reg21_out;
  wire par_done_reg21_done;
  wire par_done_reg22_in;
  wire par_done_reg22_write_en;
  wire par_done_reg22_clk;
  wire par_done_reg22_out;
  wire par_done_reg22_done;
  wire par_reset5_in;
  wire par_reset5_write_en;
  wire par_reset5_clk;
  wire par_reset5_out;
  wire par_reset5_done;
  wire par_done_reg23_in;
  wire par_done_reg23_write_en;
  wire par_done_reg23_clk;
  wire par_done_reg23_out;
  wire par_done_reg23_done;
  wire par_done_reg24_in;
  wire par_done_reg24_write_en;
  wire par_done_reg24_clk;
  wire par_done_reg24_out;
  wire par_done_reg24_done;
  wire par_done_reg25_in;
  wire par_done_reg25_write_en;
  wire par_done_reg25_clk;
  wire par_done_reg25_out;
  wire par_done_reg25_done;
  wire par_done_reg26_in;
  wire par_done_reg26_write_en;
  wire par_done_reg26_clk;
  wire par_done_reg26_out;
  wire par_done_reg26_done;
  wire par_done_reg27_in;
  wire par_done_reg27_write_en;
  wire par_done_reg27_clk;
  wire par_done_reg27_out;
  wire par_done_reg27_done;
  wire par_done_reg28_in;
  wire par_done_reg28_write_en;
  wire par_done_reg28_clk;
  wire par_done_reg28_out;
  wire par_done_reg28_done;
  wire par_done_reg29_in;
  wire par_done_reg29_write_en;
  wire par_done_reg29_clk;
  wire par_done_reg29_out;
  wire par_done_reg29_done;
  wire par_done_reg30_in;
  wire par_done_reg30_write_en;
  wire par_done_reg30_clk;
  wire par_done_reg30_out;
  wire par_done_reg30_done;
  wire par_done_reg31_in;
  wire par_done_reg31_write_en;
  wire par_done_reg31_clk;
  wire par_done_reg31_out;
  wire par_done_reg31_done;
  wire par_reset6_in;
  wire par_reset6_write_en;
  wire par_reset6_clk;
  wire par_reset6_out;
  wire par_reset6_done;
  wire par_done_reg32_in;
  wire par_done_reg32_write_en;
  wire par_done_reg32_clk;
  wire par_done_reg32_out;
  wire par_done_reg32_done;
  wire par_done_reg33_in;
  wire par_done_reg33_write_en;
  wire par_done_reg33_clk;
  wire par_done_reg33_out;
  wire par_done_reg33_done;
  wire par_done_reg34_in;
  wire par_done_reg34_write_en;
  wire par_done_reg34_clk;
  wire par_done_reg34_out;
  wire par_done_reg34_done;
  wire par_done_reg35_in;
  wire par_done_reg35_write_en;
  wire par_done_reg35_clk;
  wire par_done_reg35_out;
  wire par_done_reg35_done;
  wire par_done_reg36_in;
  wire par_done_reg36_write_en;
  wire par_done_reg36_clk;
  wire par_done_reg36_out;
  wire par_done_reg36_done;
  wire par_done_reg37_in;
  wire par_done_reg37_write_en;
  wire par_done_reg37_clk;
  wire par_done_reg37_out;
  wire par_done_reg37_done;
  wire par_done_reg38_in;
  wire par_done_reg38_write_en;
  wire par_done_reg38_clk;
  wire par_done_reg38_out;
  wire par_done_reg38_done;
  wire par_done_reg39_in;
  wire par_done_reg39_write_en;
  wire par_done_reg39_clk;
  wire par_done_reg39_out;
  wire par_done_reg39_done;
  wire par_done_reg40_in;
  wire par_done_reg40_write_en;
  wire par_done_reg40_clk;
  wire par_done_reg40_out;
  wire par_done_reg40_done;
  wire par_done_reg41_in;
  wire par_done_reg41_write_en;
  wire par_done_reg41_clk;
  wire par_done_reg41_out;
  wire par_done_reg41_done;
  wire par_done_reg42_in;
  wire par_done_reg42_write_en;
  wire par_done_reg42_clk;
  wire par_done_reg42_out;
  wire par_done_reg42_done;
  wire par_done_reg43_in;
  wire par_done_reg43_write_en;
  wire par_done_reg43_clk;
  wire par_done_reg43_out;
  wire par_done_reg43_done;
  wire par_reset7_in;
  wire par_reset7_write_en;
  wire par_reset7_clk;
  wire par_reset7_out;
  wire par_reset7_done;
  wire par_done_reg44_in;
  wire par_done_reg44_write_en;
  wire par_done_reg44_clk;
  wire par_done_reg44_out;
  wire par_done_reg44_done;
  wire par_done_reg45_in;
  wire par_done_reg45_write_en;
  wire par_done_reg45_clk;
  wire par_done_reg45_out;
  wire par_done_reg45_done;
  wire par_done_reg46_in;
  wire par_done_reg46_write_en;
  wire par_done_reg46_clk;
  wire par_done_reg46_out;
  wire par_done_reg46_done;
  wire par_done_reg47_in;
  wire par_done_reg47_write_en;
  wire par_done_reg47_clk;
  wire par_done_reg47_out;
  wire par_done_reg47_done;
  wire par_done_reg48_in;
  wire par_done_reg48_write_en;
  wire par_done_reg48_clk;
  wire par_done_reg48_out;
  wire par_done_reg48_done;
  wire par_done_reg49_in;
  wire par_done_reg49_write_en;
  wire par_done_reg49_clk;
  wire par_done_reg49_out;
  wire par_done_reg49_done;
  wire par_done_reg50_in;
  wire par_done_reg50_write_en;
  wire par_done_reg50_clk;
  wire par_done_reg50_out;
  wire par_done_reg50_done;
  wire par_done_reg51_in;
  wire par_done_reg51_write_en;
  wire par_done_reg51_clk;
  wire par_done_reg51_out;
  wire par_done_reg51_done;
  wire par_done_reg52_in;
  wire par_done_reg52_write_en;
  wire par_done_reg52_clk;
  wire par_done_reg52_out;
  wire par_done_reg52_done;
  wire par_done_reg53_in;
  wire par_done_reg53_write_en;
  wire par_done_reg53_clk;
  wire par_done_reg53_out;
  wire par_done_reg53_done;
  wire par_done_reg54_in;
  wire par_done_reg54_write_en;
  wire par_done_reg54_clk;
  wire par_done_reg54_out;
  wire par_done_reg54_done;
  wire par_done_reg55_in;
  wire par_done_reg55_write_en;
  wire par_done_reg55_clk;
  wire par_done_reg55_out;
  wire par_done_reg55_done;
  wire par_done_reg56_in;
  wire par_done_reg56_write_en;
  wire par_done_reg56_clk;
  wire par_done_reg56_out;
  wire par_done_reg56_done;
  wire par_done_reg57_in;
  wire par_done_reg57_write_en;
  wire par_done_reg57_clk;
  wire par_done_reg57_out;
  wire par_done_reg57_done;
  wire par_reset8_in;
  wire par_reset8_write_en;
  wire par_reset8_clk;
  wire par_reset8_out;
  wire par_reset8_done;
  wire par_done_reg58_in;
  wire par_done_reg58_write_en;
  wire par_done_reg58_clk;
  wire par_done_reg58_out;
  wire par_done_reg58_done;
  wire par_done_reg59_in;
  wire par_done_reg59_write_en;
  wire par_done_reg59_clk;
  wire par_done_reg59_out;
  wire par_done_reg59_done;
  wire par_done_reg60_in;
  wire par_done_reg60_write_en;
  wire par_done_reg60_clk;
  wire par_done_reg60_out;
  wire par_done_reg60_done;
  wire par_done_reg61_in;
  wire par_done_reg61_write_en;
  wire par_done_reg61_clk;
  wire par_done_reg61_out;
  wire par_done_reg61_done;
  wire par_done_reg62_in;
  wire par_done_reg62_write_en;
  wire par_done_reg62_clk;
  wire par_done_reg62_out;
  wire par_done_reg62_done;
  wire par_done_reg63_in;
  wire par_done_reg63_write_en;
  wire par_done_reg63_clk;
  wire par_done_reg63_out;
  wire par_done_reg63_done;
  wire par_done_reg64_in;
  wire par_done_reg64_write_en;
  wire par_done_reg64_clk;
  wire par_done_reg64_out;
  wire par_done_reg64_done;
  wire par_done_reg65_in;
  wire par_done_reg65_write_en;
  wire par_done_reg65_clk;
  wire par_done_reg65_out;
  wire par_done_reg65_done;
  wire par_done_reg66_in;
  wire par_done_reg66_write_en;
  wire par_done_reg66_clk;
  wire par_done_reg66_out;
  wire par_done_reg66_done;
  wire par_done_reg67_in;
  wire par_done_reg67_write_en;
  wire par_done_reg67_clk;
  wire par_done_reg67_out;
  wire par_done_reg67_done;
  wire par_done_reg68_in;
  wire par_done_reg68_write_en;
  wire par_done_reg68_clk;
  wire par_done_reg68_out;
  wire par_done_reg68_done;
  wire par_done_reg69_in;
  wire par_done_reg69_write_en;
  wire par_done_reg69_clk;
  wire par_done_reg69_out;
  wire par_done_reg69_done;
  wire par_done_reg70_in;
  wire par_done_reg70_write_en;
  wire par_done_reg70_clk;
  wire par_done_reg70_out;
  wire par_done_reg70_done;
  wire par_done_reg71_in;
  wire par_done_reg71_write_en;
  wire par_done_reg71_clk;
  wire par_done_reg71_out;
  wire par_done_reg71_done;
  wire par_done_reg72_in;
  wire par_done_reg72_write_en;
  wire par_done_reg72_clk;
  wire par_done_reg72_out;
  wire par_done_reg72_done;
  wire par_done_reg73_in;
  wire par_done_reg73_write_en;
  wire par_done_reg73_clk;
  wire par_done_reg73_out;
  wire par_done_reg73_done;
  wire par_done_reg74_in;
  wire par_done_reg74_write_en;
  wire par_done_reg74_clk;
  wire par_done_reg74_out;
  wire par_done_reg74_done;
  wire par_done_reg75_in;
  wire par_done_reg75_write_en;
  wire par_done_reg75_clk;
  wire par_done_reg75_out;
  wire par_done_reg75_done;
  wire par_done_reg76_in;
  wire par_done_reg76_write_en;
  wire par_done_reg76_clk;
  wire par_done_reg76_out;
  wire par_done_reg76_done;
  wire par_done_reg77_in;
  wire par_done_reg77_write_en;
  wire par_done_reg77_clk;
  wire par_done_reg77_out;
  wire par_done_reg77_done;
  wire par_reset9_in;
  wire par_reset9_write_en;
  wire par_reset9_clk;
  wire par_reset9_out;
  wire par_reset9_done;
  wire par_done_reg78_in;
  wire par_done_reg78_write_en;
  wire par_done_reg78_clk;
  wire par_done_reg78_out;
  wire par_done_reg78_done;
  wire par_done_reg79_in;
  wire par_done_reg79_write_en;
  wire par_done_reg79_clk;
  wire par_done_reg79_out;
  wire par_done_reg79_done;
  wire par_done_reg80_in;
  wire par_done_reg80_write_en;
  wire par_done_reg80_clk;
  wire par_done_reg80_out;
  wire par_done_reg80_done;
  wire par_done_reg81_in;
  wire par_done_reg81_write_en;
  wire par_done_reg81_clk;
  wire par_done_reg81_out;
  wire par_done_reg81_done;
  wire par_done_reg82_in;
  wire par_done_reg82_write_en;
  wire par_done_reg82_clk;
  wire par_done_reg82_out;
  wire par_done_reg82_done;
  wire par_done_reg83_in;
  wire par_done_reg83_write_en;
  wire par_done_reg83_clk;
  wire par_done_reg83_out;
  wire par_done_reg83_done;
  wire par_done_reg84_in;
  wire par_done_reg84_write_en;
  wire par_done_reg84_clk;
  wire par_done_reg84_out;
  wire par_done_reg84_done;
  wire par_done_reg85_in;
  wire par_done_reg85_write_en;
  wire par_done_reg85_clk;
  wire par_done_reg85_out;
  wire par_done_reg85_done;
  wire par_done_reg86_in;
  wire par_done_reg86_write_en;
  wire par_done_reg86_clk;
  wire par_done_reg86_out;
  wire par_done_reg86_done;
  wire par_done_reg87_in;
  wire par_done_reg87_write_en;
  wire par_done_reg87_clk;
  wire par_done_reg87_out;
  wire par_done_reg87_done;
  wire par_done_reg88_in;
  wire par_done_reg88_write_en;
  wire par_done_reg88_clk;
  wire par_done_reg88_out;
  wire par_done_reg88_done;
  wire par_done_reg89_in;
  wire par_done_reg89_write_en;
  wire par_done_reg89_clk;
  wire par_done_reg89_out;
  wire par_done_reg89_done;
  wire par_done_reg90_in;
  wire par_done_reg90_write_en;
  wire par_done_reg90_clk;
  wire par_done_reg90_out;
  wire par_done_reg90_done;
  wire par_done_reg91_in;
  wire par_done_reg91_write_en;
  wire par_done_reg91_clk;
  wire par_done_reg91_out;
  wire par_done_reg91_done;
  wire par_done_reg92_in;
  wire par_done_reg92_write_en;
  wire par_done_reg92_clk;
  wire par_done_reg92_out;
  wire par_done_reg92_done;
  wire par_done_reg93_in;
  wire par_done_reg93_write_en;
  wire par_done_reg93_clk;
  wire par_done_reg93_out;
  wire par_done_reg93_done;
  wire par_reset10_in;
  wire par_reset10_write_en;
  wire par_reset10_clk;
  wire par_reset10_out;
  wire par_reset10_done;
  wire par_done_reg94_in;
  wire par_done_reg94_write_en;
  wire par_done_reg94_clk;
  wire par_done_reg94_out;
  wire par_done_reg94_done;
  wire par_done_reg95_in;
  wire par_done_reg95_write_en;
  wire par_done_reg95_clk;
  wire par_done_reg95_out;
  wire par_done_reg95_done;
  wire par_done_reg96_in;
  wire par_done_reg96_write_en;
  wire par_done_reg96_clk;
  wire par_done_reg96_out;
  wire par_done_reg96_done;
  wire par_done_reg97_in;
  wire par_done_reg97_write_en;
  wire par_done_reg97_clk;
  wire par_done_reg97_out;
  wire par_done_reg97_done;
  wire par_done_reg98_in;
  wire par_done_reg98_write_en;
  wire par_done_reg98_clk;
  wire par_done_reg98_out;
  wire par_done_reg98_done;
  wire par_done_reg99_in;
  wire par_done_reg99_write_en;
  wire par_done_reg99_clk;
  wire par_done_reg99_out;
  wire par_done_reg99_done;
  wire par_done_reg100_in;
  wire par_done_reg100_write_en;
  wire par_done_reg100_clk;
  wire par_done_reg100_out;
  wire par_done_reg100_done;
  wire par_done_reg101_in;
  wire par_done_reg101_write_en;
  wire par_done_reg101_clk;
  wire par_done_reg101_out;
  wire par_done_reg101_done;
  wire par_done_reg102_in;
  wire par_done_reg102_write_en;
  wire par_done_reg102_clk;
  wire par_done_reg102_out;
  wire par_done_reg102_done;
  wire par_done_reg103_in;
  wire par_done_reg103_write_en;
  wire par_done_reg103_clk;
  wire par_done_reg103_out;
  wire par_done_reg103_done;
  wire par_done_reg104_in;
  wire par_done_reg104_write_en;
  wire par_done_reg104_clk;
  wire par_done_reg104_out;
  wire par_done_reg104_done;
  wire par_done_reg105_in;
  wire par_done_reg105_write_en;
  wire par_done_reg105_clk;
  wire par_done_reg105_out;
  wire par_done_reg105_done;
  wire par_done_reg106_in;
  wire par_done_reg106_write_en;
  wire par_done_reg106_clk;
  wire par_done_reg106_out;
  wire par_done_reg106_done;
  wire par_done_reg107_in;
  wire par_done_reg107_write_en;
  wire par_done_reg107_clk;
  wire par_done_reg107_out;
  wire par_done_reg107_done;
  wire par_done_reg108_in;
  wire par_done_reg108_write_en;
  wire par_done_reg108_clk;
  wire par_done_reg108_out;
  wire par_done_reg108_done;
  wire par_done_reg109_in;
  wire par_done_reg109_write_en;
  wire par_done_reg109_clk;
  wire par_done_reg109_out;
  wire par_done_reg109_done;
  wire par_done_reg110_in;
  wire par_done_reg110_write_en;
  wire par_done_reg110_clk;
  wire par_done_reg110_out;
  wire par_done_reg110_done;
  wire par_done_reg111_in;
  wire par_done_reg111_write_en;
  wire par_done_reg111_clk;
  wire par_done_reg111_out;
  wire par_done_reg111_done;
  wire par_done_reg112_in;
  wire par_done_reg112_write_en;
  wire par_done_reg112_clk;
  wire par_done_reg112_out;
  wire par_done_reg112_done;
  wire par_done_reg113_in;
  wire par_done_reg113_write_en;
  wire par_done_reg113_clk;
  wire par_done_reg113_out;
  wire par_done_reg113_done;
  wire par_done_reg114_in;
  wire par_done_reg114_write_en;
  wire par_done_reg114_clk;
  wire par_done_reg114_out;
  wire par_done_reg114_done;
  wire par_done_reg115_in;
  wire par_done_reg115_write_en;
  wire par_done_reg115_clk;
  wire par_done_reg115_out;
  wire par_done_reg115_done;
  wire par_done_reg116_in;
  wire par_done_reg116_write_en;
  wire par_done_reg116_clk;
  wire par_done_reg116_out;
  wire par_done_reg116_done;
  wire par_done_reg117_in;
  wire par_done_reg117_write_en;
  wire par_done_reg117_clk;
  wire par_done_reg117_out;
  wire par_done_reg117_done;
  wire par_reset11_in;
  wire par_reset11_write_en;
  wire par_reset11_clk;
  wire par_reset11_out;
  wire par_reset11_done;
  wire par_done_reg118_in;
  wire par_done_reg118_write_en;
  wire par_done_reg118_clk;
  wire par_done_reg118_out;
  wire par_done_reg118_done;
  wire par_done_reg119_in;
  wire par_done_reg119_write_en;
  wire par_done_reg119_clk;
  wire par_done_reg119_out;
  wire par_done_reg119_done;
  wire par_done_reg120_in;
  wire par_done_reg120_write_en;
  wire par_done_reg120_clk;
  wire par_done_reg120_out;
  wire par_done_reg120_done;
  wire par_done_reg121_in;
  wire par_done_reg121_write_en;
  wire par_done_reg121_clk;
  wire par_done_reg121_out;
  wire par_done_reg121_done;
  wire par_done_reg122_in;
  wire par_done_reg122_write_en;
  wire par_done_reg122_clk;
  wire par_done_reg122_out;
  wire par_done_reg122_done;
  wire par_done_reg123_in;
  wire par_done_reg123_write_en;
  wire par_done_reg123_clk;
  wire par_done_reg123_out;
  wire par_done_reg123_done;
  wire par_done_reg124_in;
  wire par_done_reg124_write_en;
  wire par_done_reg124_clk;
  wire par_done_reg124_out;
  wire par_done_reg124_done;
  wire par_done_reg125_in;
  wire par_done_reg125_write_en;
  wire par_done_reg125_clk;
  wire par_done_reg125_out;
  wire par_done_reg125_done;
  wire par_done_reg126_in;
  wire par_done_reg126_write_en;
  wire par_done_reg126_clk;
  wire par_done_reg126_out;
  wire par_done_reg126_done;
  wire par_done_reg127_in;
  wire par_done_reg127_write_en;
  wire par_done_reg127_clk;
  wire par_done_reg127_out;
  wire par_done_reg127_done;
  wire par_done_reg128_in;
  wire par_done_reg128_write_en;
  wire par_done_reg128_clk;
  wire par_done_reg128_out;
  wire par_done_reg128_done;
  wire par_done_reg129_in;
  wire par_done_reg129_write_en;
  wire par_done_reg129_clk;
  wire par_done_reg129_out;
  wire par_done_reg129_done;
  wire par_done_reg130_in;
  wire par_done_reg130_write_en;
  wire par_done_reg130_clk;
  wire par_done_reg130_out;
  wire par_done_reg130_done;
  wire par_done_reg131_in;
  wire par_done_reg131_write_en;
  wire par_done_reg131_clk;
  wire par_done_reg131_out;
  wire par_done_reg131_done;
  wire par_done_reg132_in;
  wire par_done_reg132_write_en;
  wire par_done_reg132_clk;
  wire par_done_reg132_out;
  wire par_done_reg132_done;
  wire par_done_reg133_in;
  wire par_done_reg133_write_en;
  wire par_done_reg133_clk;
  wire par_done_reg133_out;
  wire par_done_reg133_done;
  wire par_reset12_in;
  wire par_reset12_write_en;
  wire par_reset12_clk;
  wire par_reset12_out;
  wire par_reset12_done;
  wire par_done_reg134_in;
  wire par_done_reg134_write_en;
  wire par_done_reg134_clk;
  wire par_done_reg134_out;
  wire par_done_reg134_done;
  wire par_done_reg135_in;
  wire par_done_reg135_write_en;
  wire par_done_reg135_clk;
  wire par_done_reg135_out;
  wire par_done_reg135_done;
  wire par_done_reg136_in;
  wire par_done_reg136_write_en;
  wire par_done_reg136_clk;
  wire par_done_reg136_out;
  wire par_done_reg136_done;
  wire par_done_reg137_in;
  wire par_done_reg137_write_en;
  wire par_done_reg137_clk;
  wire par_done_reg137_out;
  wire par_done_reg137_done;
  wire par_done_reg138_in;
  wire par_done_reg138_write_en;
  wire par_done_reg138_clk;
  wire par_done_reg138_out;
  wire par_done_reg138_done;
  wire par_done_reg139_in;
  wire par_done_reg139_write_en;
  wire par_done_reg139_clk;
  wire par_done_reg139_out;
  wire par_done_reg139_done;
  wire par_done_reg140_in;
  wire par_done_reg140_write_en;
  wire par_done_reg140_clk;
  wire par_done_reg140_out;
  wire par_done_reg140_done;
  wire par_done_reg141_in;
  wire par_done_reg141_write_en;
  wire par_done_reg141_clk;
  wire par_done_reg141_out;
  wire par_done_reg141_done;
  wire par_done_reg142_in;
  wire par_done_reg142_write_en;
  wire par_done_reg142_clk;
  wire par_done_reg142_out;
  wire par_done_reg142_done;
  wire par_done_reg143_in;
  wire par_done_reg143_write_en;
  wire par_done_reg143_clk;
  wire par_done_reg143_out;
  wire par_done_reg143_done;
  wire par_done_reg144_in;
  wire par_done_reg144_write_en;
  wire par_done_reg144_clk;
  wire par_done_reg144_out;
  wire par_done_reg144_done;
  wire par_done_reg145_in;
  wire par_done_reg145_write_en;
  wire par_done_reg145_clk;
  wire par_done_reg145_out;
  wire par_done_reg145_done;
  wire par_done_reg146_in;
  wire par_done_reg146_write_en;
  wire par_done_reg146_clk;
  wire par_done_reg146_out;
  wire par_done_reg146_done;
  wire par_done_reg147_in;
  wire par_done_reg147_write_en;
  wire par_done_reg147_clk;
  wire par_done_reg147_out;
  wire par_done_reg147_done;
  wire par_done_reg148_in;
  wire par_done_reg148_write_en;
  wire par_done_reg148_clk;
  wire par_done_reg148_out;
  wire par_done_reg148_done;
  wire par_done_reg149_in;
  wire par_done_reg149_write_en;
  wire par_done_reg149_clk;
  wire par_done_reg149_out;
  wire par_done_reg149_done;
  wire par_done_reg150_in;
  wire par_done_reg150_write_en;
  wire par_done_reg150_clk;
  wire par_done_reg150_out;
  wire par_done_reg150_done;
  wire par_done_reg151_in;
  wire par_done_reg151_write_en;
  wire par_done_reg151_clk;
  wire par_done_reg151_out;
  wire par_done_reg151_done;
  wire par_done_reg152_in;
  wire par_done_reg152_write_en;
  wire par_done_reg152_clk;
  wire par_done_reg152_out;
  wire par_done_reg152_done;
  wire par_done_reg153_in;
  wire par_done_reg153_write_en;
  wire par_done_reg153_clk;
  wire par_done_reg153_out;
  wire par_done_reg153_done;
  wire par_done_reg154_in;
  wire par_done_reg154_write_en;
  wire par_done_reg154_clk;
  wire par_done_reg154_out;
  wire par_done_reg154_done;
  wire par_done_reg155_in;
  wire par_done_reg155_write_en;
  wire par_done_reg155_clk;
  wire par_done_reg155_out;
  wire par_done_reg155_done;
  wire par_done_reg156_in;
  wire par_done_reg156_write_en;
  wire par_done_reg156_clk;
  wire par_done_reg156_out;
  wire par_done_reg156_done;
  wire par_done_reg157_in;
  wire par_done_reg157_write_en;
  wire par_done_reg157_clk;
  wire par_done_reg157_out;
  wire par_done_reg157_done;
  wire par_reset13_in;
  wire par_reset13_write_en;
  wire par_reset13_clk;
  wire par_reset13_out;
  wire par_reset13_done;
  wire par_done_reg158_in;
  wire par_done_reg158_write_en;
  wire par_done_reg158_clk;
  wire par_done_reg158_out;
  wire par_done_reg158_done;
  wire par_done_reg159_in;
  wire par_done_reg159_write_en;
  wire par_done_reg159_clk;
  wire par_done_reg159_out;
  wire par_done_reg159_done;
  wire par_done_reg160_in;
  wire par_done_reg160_write_en;
  wire par_done_reg160_clk;
  wire par_done_reg160_out;
  wire par_done_reg160_done;
  wire par_done_reg161_in;
  wire par_done_reg161_write_en;
  wire par_done_reg161_clk;
  wire par_done_reg161_out;
  wire par_done_reg161_done;
  wire par_done_reg162_in;
  wire par_done_reg162_write_en;
  wire par_done_reg162_clk;
  wire par_done_reg162_out;
  wire par_done_reg162_done;
  wire par_done_reg163_in;
  wire par_done_reg163_write_en;
  wire par_done_reg163_clk;
  wire par_done_reg163_out;
  wire par_done_reg163_done;
  wire par_done_reg164_in;
  wire par_done_reg164_write_en;
  wire par_done_reg164_clk;
  wire par_done_reg164_out;
  wire par_done_reg164_done;
  wire par_done_reg165_in;
  wire par_done_reg165_write_en;
  wire par_done_reg165_clk;
  wire par_done_reg165_out;
  wire par_done_reg165_done;
  wire par_done_reg166_in;
  wire par_done_reg166_write_en;
  wire par_done_reg166_clk;
  wire par_done_reg166_out;
  wire par_done_reg166_done;
  wire par_done_reg167_in;
  wire par_done_reg167_write_en;
  wire par_done_reg167_clk;
  wire par_done_reg167_out;
  wire par_done_reg167_done;
  wire par_done_reg168_in;
  wire par_done_reg168_write_en;
  wire par_done_reg168_clk;
  wire par_done_reg168_out;
  wire par_done_reg168_done;
  wire par_done_reg169_in;
  wire par_done_reg169_write_en;
  wire par_done_reg169_clk;
  wire par_done_reg169_out;
  wire par_done_reg169_done;
  wire par_done_reg170_in;
  wire par_done_reg170_write_en;
  wire par_done_reg170_clk;
  wire par_done_reg170_out;
  wire par_done_reg170_done;
  wire par_done_reg171_in;
  wire par_done_reg171_write_en;
  wire par_done_reg171_clk;
  wire par_done_reg171_out;
  wire par_done_reg171_done;
  wire par_reset14_in;
  wire par_reset14_write_en;
  wire par_reset14_clk;
  wire par_reset14_out;
  wire par_reset14_done;
  wire par_done_reg172_in;
  wire par_done_reg172_write_en;
  wire par_done_reg172_clk;
  wire par_done_reg172_out;
  wire par_done_reg172_done;
  wire par_done_reg173_in;
  wire par_done_reg173_write_en;
  wire par_done_reg173_clk;
  wire par_done_reg173_out;
  wire par_done_reg173_done;
  wire par_done_reg174_in;
  wire par_done_reg174_write_en;
  wire par_done_reg174_clk;
  wire par_done_reg174_out;
  wire par_done_reg174_done;
  wire par_done_reg175_in;
  wire par_done_reg175_write_en;
  wire par_done_reg175_clk;
  wire par_done_reg175_out;
  wire par_done_reg175_done;
  wire par_done_reg176_in;
  wire par_done_reg176_write_en;
  wire par_done_reg176_clk;
  wire par_done_reg176_out;
  wire par_done_reg176_done;
  wire par_done_reg177_in;
  wire par_done_reg177_write_en;
  wire par_done_reg177_clk;
  wire par_done_reg177_out;
  wire par_done_reg177_done;
  wire par_done_reg178_in;
  wire par_done_reg178_write_en;
  wire par_done_reg178_clk;
  wire par_done_reg178_out;
  wire par_done_reg178_done;
  wire par_done_reg179_in;
  wire par_done_reg179_write_en;
  wire par_done_reg179_clk;
  wire par_done_reg179_out;
  wire par_done_reg179_done;
  wire par_done_reg180_in;
  wire par_done_reg180_write_en;
  wire par_done_reg180_clk;
  wire par_done_reg180_out;
  wire par_done_reg180_done;
  wire par_done_reg181_in;
  wire par_done_reg181_write_en;
  wire par_done_reg181_clk;
  wire par_done_reg181_out;
  wire par_done_reg181_done;
  wire par_done_reg182_in;
  wire par_done_reg182_write_en;
  wire par_done_reg182_clk;
  wire par_done_reg182_out;
  wire par_done_reg182_done;
  wire par_done_reg183_in;
  wire par_done_reg183_write_en;
  wire par_done_reg183_clk;
  wire par_done_reg183_out;
  wire par_done_reg183_done;
  wire par_done_reg184_in;
  wire par_done_reg184_write_en;
  wire par_done_reg184_clk;
  wire par_done_reg184_out;
  wire par_done_reg184_done;
  wire par_done_reg185_in;
  wire par_done_reg185_write_en;
  wire par_done_reg185_clk;
  wire par_done_reg185_out;
  wire par_done_reg185_done;
  wire par_done_reg186_in;
  wire par_done_reg186_write_en;
  wire par_done_reg186_clk;
  wire par_done_reg186_out;
  wire par_done_reg186_done;
  wire par_done_reg187_in;
  wire par_done_reg187_write_en;
  wire par_done_reg187_clk;
  wire par_done_reg187_out;
  wire par_done_reg187_done;
  wire par_done_reg188_in;
  wire par_done_reg188_write_en;
  wire par_done_reg188_clk;
  wire par_done_reg188_out;
  wire par_done_reg188_done;
  wire par_done_reg189_in;
  wire par_done_reg189_write_en;
  wire par_done_reg189_clk;
  wire par_done_reg189_out;
  wire par_done_reg189_done;
  wire par_done_reg190_in;
  wire par_done_reg190_write_en;
  wire par_done_reg190_clk;
  wire par_done_reg190_out;
  wire par_done_reg190_done;
  wire par_done_reg191_in;
  wire par_done_reg191_write_en;
  wire par_done_reg191_clk;
  wire par_done_reg191_out;
  wire par_done_reg191_done;
  wire par_reset15_in;
  wire par_reset15_write_en;
  wire par_reset15_clk;
  wire par_reset15_out;
  wire par_reset15_done;
  wire par_done_reg192_in;
  wire par_done_reg192_write_en;
  wire par_done_reg192_clk;
  wire par_done_reg192_out;
  wire par_done_reg192_done;
  wire par_done_reg193_in;
  wire par_done_reg193_write_en;
  wire par_done_reg193_clk;
  wire par_done_reg193_out;
  wire par_done_reg193_done;
  wire par_done_reg194_in;
  wire par_done_reg194_write_en;
  wire par_done_reg194_clk;
  wire par_done_reg194_out;
  wire par_done_reg194_done;
  wire par_done_reg195_in;
  wire par_done_reg195_write_en;
  wire par_done_reg195_clk;
  wire par_done_reg195_out;
  wire par_done_reg195_done;
  wire par_done_reg196_in;
  wire par_done_reg196_write_en;
  wire par_done_reg196_clk;
  wire par_done_reg196_out;
  wire par_done_reg196_done;
  wire par_done_reg197_in;
  wire par_done_reg197_write_en;
  wire par_done_reg197_clk;
  wire par_done_reg197_out;
  wire par_done_reg197_done;
  wire par_done_reg198_in;
  wire par_done_reg198_write_en;
  wire par_done_reg198_clk;
  wire par_done_reg198_out;
  wire par_done_reg198_done;
  wire par_done_reg199_in;
  wire par_done_reg199_write_en;
  wire par_done_reg199_clk;
  wire par_done_reg199_out;
  wire par_done_reg199_done;
  wire par_done_reg200_in;
  wire par_done_reg200_write_en;
  wire par_done_reg200_clk;
  wire par_done_reg200_out;
  wire par_done_reg200_done;
  wire par_done_reg201_in;
  wire par_done_reg201_write_en;
  wire par_done_reg201_clk;
  wire par_done_reg201_out;
  wire par_done_reg201_done;
  wire par_reset16_in;
  wire par_reset16_write_en;
  wire par_reset16_clk;
  wire par_reset16_out;
  wire par_reset16_done;
  wire par_done_reg202_in;
  wire par_done_reg202_write_en;
  wire par_done_reg202_clk;
  wire par_done_reg202_out;
  wire par_done_reg202_done;
  wire par_done_reg203_in;
  wire par_done_reg203_write_en;
  wire par_done_reg203_clk;
  wire par_done_reg203_out;
  wire par_done_reg203_done;
  wire par_done_reg204_in;
  wire par_done_reg204_write_en;
  wire par_done_reg204_clk;
  wire par_done_reg204_out;
  wire par_done_reg204_done;
  wire par_done_reg205_in;
  wire par_done_reg205_write_en;
  wire par_done_reg205_clk;
  wire par_done_reg205_out;
  wire par_done_reg205_done;
  wire par_done_reg206_in;
  wire par_done_reg206_write_en;
  wire par_done_reg206_clk;
  wire par_done_reg206_out;
  wire par_done_reg206_done;
  wire par_done_reg207_in;
  wire par_done_reg207_write_en;
  wire par_done_reg207_clk;
  wire par_done_reg207_out;
  wire par_done_reg207_done;
  wire par_done_reg208_in;
  wire par_done_reg208_write_en;
  wire par_done_reg208_clk;
  wire par_done_reg208_out;
  wire par_done_reg208_done;
  wire par_done_reg209_in;
  wire par_done_reg209_write_en;
  wire par_done_reg209_clk;
  wire par_done_reg209_out;
  wire par_done_reg209_done;
  wire par_done_reg210_in;
  wire par_done_reg210_write_en;
  wire par_done_reg210_clk;
  wire par_done_reg210_out;
  wire par_done_reg210_done;
  wire par_done_reg211_in;
  wire par_done_reg211_write_en;
  wire par_done_reg211_clk;
  wire par_done_reg211_out;
  wire par_done_reg211_done;
  wire par_done_reg212_in;
  wire par_done_reg212_write_en;
  wire par_done_reg212_clk;
  wire par_done_reg212_out;
  wire par_done_reg212_done;
  wire par_done_reg213_in;
  wire par_done_reg213_write_en;
  wire par_done_reg213_clk;
  wire par_done_reg213_out;
  wire par_done_reg213_done;
  wire par_reset17_in;
  wire par_reset17_write_en;
  wire par_reset17_clk;
  wire par_reset17_out;
  wire par_reset17_done;
  wire par_done_reg214_in;
  wire par_done_reg214_write_en;
  wire par_done_reg214_clk;
  wire par_done_reg214_out;
  wire par_done_reg214_done;
  wire par_done_reg215_in;
  wire par_done_reg215_write_en;
  wire par_done_reg215_clk;
  wire par_done_reg215_out;
  wire par_done_reg215_done;
  wire par_done_reg216_in;
  wire par_done_reg216_write_en;
  wire par_done_reg216_clk;
  wire par_done_reg216_out;
  wire par_done_reg216_done;
  wire par_done_reg217_in;
  wire par_done_reg217_write_en;
  wire par_done_reg217_clk;
  wire par_done_reg217_out;
  wire par_done_reg217_done;
  wire par_done_reg218_in;
  wire par_done_reg218_write_en;
  wire par_done_reg218_clk;
  wire par_done_reg218_out;
  wire par_done_reg218_done;
  wire par_done_reg219_in;
  wire par_done_reg219_write_en;
  wire par_done_reg219_clk;
  wire par_done_reg219_out;
  wire par_done_reg219_done;
  wire par_reset18_in;
  wire par_reset18_write_en;
  wire par_reset18_clk;
  wire par_reset18_out;
  wire par_reset18_done;
  wire par_done_reg220_in;
  wire par_done_reg220_write_en;
  wire par_done_reg220_clk;
  wire par_done_reg220_out;
  wire par_done_reg220_done;
  wire par_done_reg221_in;
  wire par_done_reg221_write_en;
  wire par_done_reg221_clk;
  wire par_done_reg221_out;
  wire par_done_reg221_done;
  wire par_done_reg222_in;
  wire par_done_reg222_write_en;
  wire par_done_reg222_clk;
  wire par_done_reg222_out;
  wire par_done_reg222_done;
  wire par_done_reg223_in;
  wire par_done_reg223_write_en;
  wire par_done_reg223_clk;
  wire par_done_reg223_out;
  wire par_done_reg223_done;
  wire par_done_reg224_in;
  wire par_done_reg224_write_en;
  wire par_done_reg224_clk;
  wire par_done_reg224_out;
  wire par_done_reg224_done;
  wire par_done_reg225_in;
  wire par_done_reg225_write_en;
  wire par_done_reg225_clk;
  wire par_done_reg225_out;
  wire par_done_reg225_done;
  wire par_reset19_in;
  wire par_reset19_write_en;
  wire par_reset19_clk;
  wire par_reset19_out;
  wire par_reset19_done;
  wire par_done_reg226_in;
  wire par_done_reg226_write_en;
  wire par_done_reg226_clk;
  wire par_done_reg226_out;
  wire par_done_reg226_done;
  wire par_done_reg227_in;
  wire par_done_reg227_write_en;
  wire par_done_reg227_clk;
  wire par_done_reg227_out;
  wire par_done_reg227_done;
  wire par_done_reg228_in;
  wire par_done_reg228_write_en;
  wire par_done_reg228_clk;
  wire par_done_reg228_out;
  wire par_done_reg228_done;
  wire par_reset20_in;
  wire par_reset20_write_en;
  wire par_reset20_clk;
  wire par_reset20_out;
  wire par_reset20_done;
  wire par_done_reg229_in;
  wire par_done_reg229_write_en;
  wire par_done_reg229_clk;
  wire par_done_reg229_out;
  wire par_done_reg229_done;
  wire par_done_reg230_in;
  wire par_done_reg230_write_en;
  wire par_done_reg230_clk;
  wire par_done_reg230_out;
  wire par_done_reg230_done;
  wire par_reset21_in;
  wire par_reset21_write_en;
  wire par_reset21_clk;
  wire par_reset21_out;
  wire par_reset21_done;
  wire par_done_reg231_in;
  wire par_done_reg231_write_en;
  wire par_done_reg231_clk;
  wire par_done_reg231_out;
  wire par_done_reg231_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_reg #(32) left_33_read (
      .in(left_33_read_in),
      .write_en(left_33_read_write_en),
      .clk(clk),
      .out(left_33_read_out),
      .done(left_33_read_done)
  );
  
  std_reg #(32) top_33_read (
      .in(top_33_read_in),
      .write_en(top_33_read_write_en),
      .clk(clk),
      .out(top_33_read_out),
      .done(top_33_read_done)
  );
  
  mac_pe #() pe_33 (
      .top(pe_33_top),
      .left(pe_33_left),
      .go(pe_33_go),
      .clk(clk),
      .down(pe_33_down),
      .right(pe_33_right),
      .out(pe_33_out),
      .done(pe_33_done)
  );
  
  std_reg #(32) right_32_write (
      .in(right_32_write_in),
      .write_en(right_32_write_write_en),
      .clk(clk),
      .out(right_32_write_out),
      .done(right_32_write_done)
  );
  
  std_reg #(32) left_32_read (
      .in(left_32_read_in),
      .write_en(left_32_read_write_en),
      .clk(clk),
      .out(left_32_read_out),
      .done(left_32_read_done)
  );
  
  std_reg #(32) top_32_read (
      .in(top_32_read_in),
      .write_en(top_32_read_write_en),
      .clk(clk),
      .out(top_32_read_out),
      .done(top_32_read_done)
  );
  
  mac_pe #() pe_32 (
      .top(pe_32_top),
      .left(pe_32_left),
      .go(pe_32_go),
      .clk(clk),
      .down(pe_32_down),
      .right(pe_32_right),
      .out(pe_32_out),
      .done(pe_32_done)
  );
  
  std_reg #(32) right_31_write (
      .in(right_31_write_in),
      .write_en(right_31_write_write_en),
      .clk(clk),
      .out(right_31_write_out),
      .done(right_31_write_done)
  );
  
  std_reg #(32) left_31_read (
      .in(left_31_read_in),
      .write_en(left_31_read_write_en),
      .clk(clk),
      .out(left_31_read_out),
      .done(left_31_read_done)
  );
  
  std_reg #(32) top_31_read (
      .in(top_31_read_in),
      .write_en(top_31_read_write_en),
      .clk(clk),
      .out(top_31_read_out),
      .done(top_31_read_done)
  );
  
  mac_pe #() pe_31 (
      .top(pe_31_top),
      .left(pe_31_left),
      .go(pe_31_go),
      .clk(clk),
      .down(pe_31_down),
      .right(pe_31_right),
      .out(pe_31_out),
      .done(pe_31_done)
  );
  
  std_reg #(32) right_30_write (
      .in(right_30_write_in),
      .write_en(right_30_write_write_en),
      .clk(clk),
      .out(right_30_write_out),
      .done(right_30_write_done)
  );
  
  std_reg #(32) left_30_read (
      .in(left_30_read_in),
      .write_en(left_30_read_write_en),
      .clk(clk),
      .out(left_30_read_out),
      .done(left_30_read_done)
  );
  
  std_reg #(32) top_30_read (
      .in(top_30_read_in),
      .write_en(top_30_read_write_en),
      .clk(clk),
      .out(top_30_read_out),
      .done(top_30_read_done)
  );
  
  mac_pe #() pe_30 (
      .top(pe_30_top),
      .left(pe_30_left),
      .go(pe_30_go),
      .clk(clk),
      .down(pe_30_down),
      .right(pe_30_right),
      .out(pe_30_out),
      .done(pe_30_done)
  );
  
  std_reg #(32) down_23_write (
      .in(down_23_write_in),
      .write_en(down_23_write_write_en),
      .clk(clk),
      .out(down_23_write_out),
      .done(down_23_write_done)
  );
  
  std_reg #(32) left_23_read (
      .in(left_23_read_in),
      .write_en(left_23_read_write_en),
      .clk(clk),
      .out(left_23_read_out),
      .done(left_23_read_done)
  );
  
  std_reg #(32) top_23_read (
      .in(top_23_read_in),
      .write_en(top_23_read_write_en),
      .clk(clk),
      .out(top_23_read_out),
      .done(top_23_read_done)
  );
  
  mac_pe #() pe_23 (
      .top(pe_23_top),
      .left(pe_23_left),
      .go(pe_23_go),
      .clk(clk),
      .down(pe_23_down),
      .right(pe_23_right),
      .out(pe_23_out),
      .done(pe_23_done)
  );
  
  std_reg #(32) down_22_write (
      .in(down_22_write_in),
      .write_en(down_22_write_write_en),
      .clk(clk),
      .out(down_22_write_out),
      .done(down_22_write_done)
  );
  
  std_reg #(32) right_22_write (
      .in(right_22_write_in),
      .write_en(right_22_write_write_en),
      .clk(clk),
      .out(right_22_write_out),
      .done(right_22_write_done)
  );
  
  std_reg #(32) left_22_read (
      .in(left_22_read_in),
      .write_en(left_22_read_write_en),
      .clk(clk),
      .out(left_22_read_out),
      .done(left_22_read_done)
  );
  
  std_reg #(32) top_22_read (
      .in(top_22_read_in),
      .write_en(top_22_read_write_en),
      .clk(clk),
      .out(top_22_read_out),
      .done(top_22_read_done)
  );
  
  mac_pe #() pe_22 (
      .top(pe_22_top),
      .left(pe_22_left),
      .go(pe_22_go),
      .clk(clk),
      .down(pe_22_down),
      .right(pe_22_right),
      .out(pe_22_out),
      .done(pe_22_done)
  );
  
  std_reg #(32) down_21_write (
      .in(down_21_write_in),
      .write_en(down_21_write_write_en),
      .clk(clk),
      .out(down_21_write_out),
      .done(down_21_write_done)
  );
  
  std_reg #(32) right_21_write (
      .in(right_21_write_in),
      .write_en(right_21_write_write_en),
      .clk(clk),
      .out(right_21_write_out),
      .done(right_21_write_done)
  );
  
  std_reg #(32) left_21_read (
      .in(left_21_read_in),
      .write_en(left_21_read_write_en),
      .clk(clk),
      .out(left_21_read_out),
      .done(left_21_read_done)
  );
  
  std_reg #(32) top_21_read (
      .in(top_21_read_in),
      .write_en(top_21_read_write_en),
      .clk(clk),
      .out(top_21_read_out),
      .done(top_21_read_done)
  );
  
  mac_pe #() pe_21 (
      .top(pe_21_top),
      .left(pe_21_left),
      .go(pe_21_go),
      .clk(clk),
      .down(pe_21_down),
      .right(pe_21_right),
      .out(pe_21_out),
      .done(pe_21_done)
  );
  
  std_reg #(32) down_20_write (
      .in(down_20_write_in),
      .write_en(down_20_write_write_en),
      .clk(clk),
      .out(down_20_write_out),
      .done(down_20_write_done)
  );
  
  std_reg #(32) right_20_write (
      .in(right_20_write_in),
      .write_en(right_20_write_write_en),
      .clk(clk),
      .out(right_20_write_out),
      .done(right_20_write_done)
  );
  
  std_reg #(32) left_20_read (
      .in(left_20_read_in),
      .write_en(left_20_read_write_en),
      .clk(clk),
      .out(left_20_read_out),
      .done(left_20_read_done)
  );
  
  std_reg #(32) top_20_read (
      .in(top_20_read_in),
      .write_en(top_20_read_write_en),
      .clk(clk),
      .out(top_20_read_out),
      .done(top_20_read_done)
  );
  
  mac_pe #() pe_20 (
      .top(pe_20_top),
      .left(pe_20_left),
      .go(pe_20_go),
      .clk(clk),
      .down(pe_20_down),
      .right(pe_20_right),
      .out(pe_20_out),
      .done(pe_20_done)
  );
  
  std_reg #(32) down_13_write (
      .in(down_13_write_in),
      .write_en(down_13_write_write_en),
      .clk(clk),
      .out(down_13_write_out),
      .done(down_13_write_done)
  );
  
  std_reg #(32) left_13_read (
      .in(left_13_read_in),
      .write_en(left_13_read_write_en),
      .clk(clk),
      .out(left_13_read_out),
      .done(left_13_read_done)
  );
  
  std_reg #(32) top_13_read (
      .in(top_13_read_in),
      .write_en(top_13_read_write_en),
      .clk(clk),
      .out(top_13_read_out),
      .done(top_13_read_done)
  );
  
  mac_pe #() pe_13 (
      .top(pe_13_top),
      .left(pe_13_left),
      .go(pe_13_go),
      .clk(clk),
      .down(pe_13_down),
      .right(pe_13_right),
      .out(pe_13_out),
      .done(pe_13_done)
  );
  
  std_reg #(32) down_12_write (
      .in(down_12_write_in),
      .write_en(down_12_write_write_en),
      .clk(clk),
      .out(down_12_write_out),
      .done(down_12_write_done)
  );
  
  std_reg #(32) right_12_write (
      .in(right_12_write_in),
      .write_en(right_12_write_write_en),
      .clk(clk),
      .out(right_12_write_out),
      .done(right_12_write_done)
  );
  
  std_reg #(32) left_12_read (
      .in(left_12_read_in),
      .write_en(left_12_read_write_en),
      .clk(clk),
      .out(left_12_read_out),
      .done(left_12_read_done)
  );
  
  std_reg #(32) top_12_read (
      .in(top_12_read_in),
      .write_en(top_12_read_write_en),
      .clk(clk),
      .out(top_12_read_out),
      .done(top_12_read_done)
  );
  
  mac_pe #() pe_12 (
      .top(pe_12_top),
      .left(pe_12_left),
      .go(pe_12_go),
      .clk(clk),
      .down(pe_12_down),
      .right(pe_12_right),
      .out(pe_12_out),
      .done(pe_12_done)
  );
  
  std_reg #(32) down_11_write (
      .in(down_11_write_in),
      .write_en(down_11_write_write_en),
      .clk(clk),
      .out(down_11_write_out),
      .done(down_11_write_done)
  );
  
  std_reg #(32) right_11_write (
      .in(right_11_write_in),
      .write_en(right_11_write_write_en),
      .clk(clk),
      .out(right_11_write_out),
      .done(right_11_write_done)
  );
  
  std_reg #(32) left_11_read (
      .in(left_11_read_in),
      .write_en(left_11_read_write_en),
      .clk(clk),
      .out(left_11_read_out),
      .done(left_11_read_done)
  );
  
  std_reg #(32) top_11_read (
      .in(top_11_read_in),
      .write_en(top_11_read_write_en),
      .clk(clk),
      .out(top_11_read_out),
      .done(top_11_read_done)
  );
  
  mac_pe #() pe_11 (
      .top(pe_11_top),
      .left(pe_11_left),
      .go(pe_11_go),
      .clk(clk),
      .down(pe_11_down),
      .right(pe_11_right),
      .out(pe_11_out),
      .done(pe_11_done)
  );
  
  std_reg #(32) down_10_write (
      .in(down_10_write_in),
      .write_en(down_10_write_write_en),
      .clk(clk),
      .out(down_10_write_out),
      .done(down_10_write_done)
  );
  
  std_reg #(32) right_10_write (
      .in(right_10_write_in),
      .write_en(right_10_write_write_en),
      .clk(clk),
      .out(right_10_write_out),
      .done(right_10_write_done)
  );
  
  std_reg #(32) left_10_read (
      .in(left_10_read_in),
      .write_en(left_10_read_write_en),
      .clk(clk),
      .out(left_10_read_out),
      .done(left_10_read_done)
  );
  
  std_reg #(32) top_10_read (
      .in(top_10_read_in),
      .write_en(top_10_read_write_en),
      .clk(clk),
      .out(top_10_read_out),
      .done(top_10_read_done)
  );
  
  mac_pe #() pe_10 (
      .top(pe_10_top),
      .left(pe_10_left),
      .go(pe_10_go),
      .clk(clk),
      .down(pe_10_down),
      .right(pe_10_right),
      .out(pe_10_out),
      .done(pe_10_done)
  );
  
  std_reg #(32) down_03_write (
      .in(down_03_write_in),
      .write_en(down_03_write_write_en),
      .clk(clk),
      .out(down_03_write_out),
      .done(down_03_write_done)
  );
  
  std_reg #(32) left_03_read (
      .in(left_03_read_in),
      .write_en(left_03_read_write_en),
      .clk(clk),
      .out(left_03_read_out),
      .done(left_03_read_done)
  );
  
  std_reg #(32) top_03_read (
      .in(top_03_read_in),
      .write_en(top_03_read_write_en),
      .clk(clk),
      .out(top_03_read_out),
      .done(top_03_read_done)
  );
  
  mac_pe #() pe_03 (
      .top(pe_03_top),
      .left(pe_03_left),
      .go(pe_03_go),
      .clk(clk),
      .down(pe_03_down),
      .right(pe_03_right),
      .out(pe_03_out),
      .done(pe_03_done)
  );
  
  std_reg #(32) down_02_write (
      .in(down_02_write_in),
      .write_en(down_02_write_write_en),
      .clk(clk),
      .out(down_02_write_out),
      .done(down_02_write_done)
  );
  
  std_reg #(32) right_02_write (
      .in(right_02_write_in),
      .write_en(right_02_write_write_en),
      .clk(clk),
      .out(right_02_write_out),
      .done(right_02_write_done)
  );
  
  std_reg #(32) left_02_read (
      .in(left_02_read_in),
      .write_en(left_02_read_write_en),
      .clk(clk),
      .out(left_02_read_out),
      .done(left_02_read_done)
  );
  
  std_reg #(32) top_02_read (
      .in(top_02_read_in),
      .write_en(top_02_read_write_en),
      .clk(clk),
      .out(top_02_read_out),
      .done(top_02_read_done)
  );
  
  mac_pe #() pe_02 (
      .top(pe_02_top),
      .left(pe_02_left),
      .go(pe_02_go),
      .clk(clk),
      .down(pe_02_down),
      .right(pe_02_right),
      .out(pe_02_out),
      .done(pe_02_done)
  );
  
  std_reg #(32) down_01_write (
      .in(down_01_write_in),
      .write_en(down_01_write_write_en),
      .clk(clk),
      .out(down_01_write_out),
      .done(down_01_write_done)
  );
  
  std_reg #(32) right_01_write (
      .in(right_01_write_in),
      .write_en(right_01_write_write_en),
      .clk(clk),
      .out(right_01_write_out),
      .done(right_01_write_done)
  );
  
  std_reg #(32) left_01_read (
      .in(left_01_read_in),
      .write_en(left_01_read_write_en),
      .clk(clk),
      .out(left_01_read_out),
      .done(left_01_read_done)
  );
  
  std_reg #(32) top_01_read (
      .in(top_01_read_in),
      .write_en(top_01_read_write_en),
      .clk(clk),
      .out(top_01_read_out),
      .done(top_01_read_done)
  );
  
  mac_pe #() pe_01 (
      .top(pe_01_top),
      .left(pe_01_left),
      .go(pe_01_go),
      .clk(clk),
      .down(pe_01_down),
      .right(pe_01_right),
      .out(pe_01_out),
      .done(pe_01_done)
  );
  
  std_reg #(32) down_00_write (
      .in(down_00_write_in),
      .write_en(down_00_write_write_en),
      .clk(clk),
      .out(down_00_write_out),
      .done(down_00_write_done)
  );
  
  std_reg #(32) right_00_write (
      .in(right_00_write_in),
      .write_en(right_00_write_write_en),
      .clk(clk),
      .out(right_00_write_out),
      .done(right_00_write_done)
  );
  
  std_reg #(32) left_00_read (
      .in(left_00_read_in),
      .write_en(left_00_read_write_en),
      .clk(clk),
      .out(left_00_read_out),
      .done(left_00_read_done)
  );
  
  std_reg #(32) top_00_read (
      .in(top_00_read_in),
      .write_en(top_00_read_write_en),
      .clk(clk),
      .out(top_00_read_out),
      .done(top_00_read_done)
  );
  
  mac_pe #() pe_00 (
      .top(pe_00_top),
      .left(pe_00_left),
      .go(pe_00_go),
      .clk(clk),
      .down(pe_00_down),
      .right(pe_00_right),
      .out(pe_00_out),
      .done(pe_00_done)
  );
  
  std_mem_d1 #(32, 4, 3) l3 (
      .addr0(l3_addr0),
      .write_data(l3_write_data),
      .write_en(l3_write_en),
      .clk(clk),
      .read_data(l3_read_data),
      .done(l3_done)
  );
  
  std_add #(3) l3_add (
      .left(l3_add_left),
      .right(l3_add_right),
      .out(l3_add_out)
  );
  
  std_reg #(3) l3_idx (
      .in(l3_idx_in),
      .write_en(l3_idx_write_en),
      .clk(clk),
      .out(l3_idx_out),
      .done(l3_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) l2 (
      .addr0(l2_addr0),
      .write_data(l2_write_data),
      .write_en(l2_write_en),
      .clk(clk),
      .read_data(l2_read_data),
      .done(l2_done)
  );
  
  std_add #(3) l2_add (
      .left(l2_add_left),
      .right(l2_add_right),
      .out(l2_add_out)
  );
  
  std_reg #(3) l2_idx (
      .in(l2_idx_in),
      .write_en(l2_idx_write_en),
      .clk(clk),
      .out(l2_idx_out),
      .done(l2_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) l1 (
      .addr0(l1_addr0),
      .write_data(l1_write_data),
      .write_en(l1_write_en),
      .clk(clk),
      .read_data(l1_read_data),
      .done(l1_done)
  );
  
  std_add #(3) l1_add (
      .left(l1_add_left),
      .right(l1_add_right),
      .out(l1_add_out)
  );
  
  std_reg #(3) l1_idx (
      .in(l1_idx_in),
      .write_en(l1_idx_write_en),
      .clk(clk),
      .out(l1_idx_out),
      .done(l1_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) l0 (
      .addr0(l0_addr0),
      .write_data(l0_write_data),
      .write_en(l0_write_en),
      .clk(clk),
      .read_data(l0_read_data),
      .done(l0_done)
  );
  
  std_add #(3) l0_add (
      .left(l0_add_left),
      .right(l0_add_right),
      .out(l0_add_out)
  );
  
  std_reg #(3) l0_idx (
      .in(l0_idx_in),
      .write_en(l0_idx_write_en),
      .clk(clk),
      .out(l0_idx_out),
      .done(l0_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) t3 (
      .addr0(t3_addr0),
      .write_data(t3_write_data),
      .write_en(t3_write_en),
      .clk(clk),
      .read_data(t3_read_data),
      .done(t3_done)
  );
  
  std_add #(3) t3_add (
      .left(t3_add_left),
      .right(t3_add_right),
      .out(t3_add_out)
  );
  
  std_reg #(3) t3_idx (
      .in(t3_idx_in),
      .write_en(t3_idx_write_en),
      .clk(clk),
      .out(t3_idx_out),
      .done(t3_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) t2 (
      .addr0(t2_addr0),
      .write_data(t2_write_data),
      .write_en(t2_write_en),
      .clk(clk),
      .read_data(t2_read_data),
      .done(t2_done)
  );
  
  std_add #(3) t2_add (
      .left(t2_add_left),
      .right(t2_add_right),
      .out(t2_add_out)
  );
  
  std_reg #(3) t2_idx (
      .in(t2_idx_in),
      .write_en(t2_idx_write_en),
      .clk(clk),
      .out(t2_idx_out),
      .done(t2_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) t1 (
      .addr0(t1_addr0),
      .write_data(t1_write_data),
      .write_en(t1_write_en),
      .clk(clk),
      .read_data(t1_read_data),
      .done(t1_done)
  );
  
  std_add #(3) t1_add (
      .left(t1_add_left),
      .right(t1_add_right),
      .out(t1_add_out)
  );
  
  std_reg #(3) t1_idx (
      .in(t1_idx_in),
      .write_en(t1_idx_write_en),
      .clk(clk),
      .out(t1_idx_out),
      .done(t1_idx_done)
  );
  
  std_mem_d1 #(32, 4, 3) t0 (
      .addr0(t0_addr0),
      .write_data(t0_write_data),
      .write_en(t0_write_en),
      .clk(clk),
      .read_data(t0_read_data),
      .done(t0_done)
  );
  
  std_add #(3) t0_add (
      .left(t0_add_left),
      .right(t0_add_right),
      .out(t0_add_out)
  );
  
  std_reg #(3) t0_idx (
      .in(t0_idx_in),
      .write_en(t0_idx_write_en),
      .clk(clk),
      .out(t0_idx_out),
      .done(t0_idx_done)
  );
  
  std_reg #(1) par_reset0 (
      .in(par_reset0_in),
      .write_en(par_reset0_write_en),
      .clk(clk),
      .out(par_reset0_out),
      .done(par_reset0_done)
  );
  
  std_reg #(1) par_done_reg0 (
      .in(par_done_reg0_in),
      .write_en(par_done_reg0_write_en),
      .clk(clk),
      .out(par_done_reg0_out),
      .done(par_done_reg0_done)
  );
  
  std_reg #(1) par_done_reg1 (
      .in(par_done_reg1_in),
      .write_en(par_done_reg1_write_en),
      .clk(clk),
      .out(par_done_reg1_out),
      .done(par_done_reg1_done)
  );
  
  std_reg #(1) par_done_reg2 (
      .in(par_done_reg2_in),
      .write_en(par_done_reg2_write_en),
      .clk(clk),
      .out(par_done_reg2_out),
      .done(par_done_reg2_done)
  );
  
  std_reg #(1) par_done_reg3 (
      .in(par_done_reg3_in),
      .write_en(par_done_reg3_write_en),
      .clk(clk),
      .out(par_done_reg3_out),
      .done(par_done_reg3_done)
  );
  
  std_reg #(1) par_done_reg4 (
      .in(par_done_reg4_in),
      .write_en(par_done_reg4_write_en),
      .clk(clk),
      .out(par_done_reg4_out),
      .done(par_done_reg4_done)
  );
  
  std_reg #(1) par_done_reg5 (
      .in(par_done_reg5_in),
      .write_en(par_done_reg5_write_en),
      .clk(clk),
      .out(par_done_reg5_out),
      .done(par_done_reg5_done)
  );
  
  std_reg #(1) par_done_reg6 (
      .in(par_done_reg6_in),
      .write_en(par_done_reg6_write_en),
      .clk(clk),
      .out(par_done_reg6_out),
      .done(par_done_reg6_done)
  );
  
  std_reg #(1) par_done_reg7 (
      .in(par_done_reg7_in),
      .write_en(par_done_reg7_write_en),
      .clk(clk),
      .out(par_done_reg7_out),
      .done(par_done_reg7_done)
  );
  
  std_reg #(1) par_reset1 (
      .in(par_reset1_in),
      .write_en(par_reset1_write_en),
      .clk(clk),
      .out(par_reset1_out),
      .done(par_reset1_done)
  );
  
  std_reg #(1) par_done_reg8 (
      .in(par_done_reg8_in),
      .write_en(par_done_reg8_write_en),
      .clk(clk),
      .out(par_done_reg8_out),
      .done(par_done_reg8_done)
  );
  
  std_reg #(1) par_done_reg9 (
      .in(par_done_reg9_in),
      .write_en(par_done_reg9_write_en),
      .clk(clk),
      .out(par_done_reg9_out),
      .done(par_done_reg9_done)
  );
  
  std_reg #(1) par_reset2 (
      .in(par_reset2_in),
      .write_en(par_reset2_write_en),
      .clk(clk),
      .out(par_reset2_out),
      .done(par_reset2_done)
  );
  
  std_reg #(1) par_done_reg10 (
      .in(par_done_reg10_in),
      .write_en(par_done_reg10_write_en),
      .clk(clk),
      .out(par_done_reg10_out),
      .done(par_done_reg10_done)
  );
  
  std_reg #(1) par_done_reg11 (
      .in(par_done_reg11_in),
      .write_en(par_done_reg11_write_en),
      .clk(clk),
      .out(par_done_reg11_out),
      .done(par_done_reg11_done)
  );
  
  std_reg #(1) par_reset3 (
      .in(par_reset3_in),
      .write_en(par_reset3_write_en),
      .clk(clk),
      .out(par_reset3_out),
      .done(par_reset3_done)
  );
  
  std_reg #(1) par_done_reg12 (
      .in(par_done_reg12_in),
      .write_en(par_done_reg12_write_en),
      .clk(clk),
      .out(par_done_reg12_out),
      .done(par_done_reg12_done)
  );
  
  std_reg #(1) par_done_reg13 (
      .in(par_done_reg13_in),
      .write_en(par_done_reg13_write_en),
      .clk(clk),
      .out(par_done_reg13_out),
      .done(par_done_reg13_done)
  );
  
  std_reg #(1) par_done_reg14 (
      .in(par_done_reg14_in),
      .write_en(par_done_reg14_write_en),
      .clk(clk),
      .out(par_done_reg14_out),
      .done(par_done_reg14_done)
  );
  
  std_reg #(1) par_done_reg15 (
      .in(par_done_reg15_in),
      .write_en(par_done_reg15_write_en),
      .clk(clk),
      .out(par_done_reg15_out),
      .done(par_done_reg15_done)
  );
  
  std_reg #(1) par_done_reg16 (
      .in(par_done_reg16_in),
      .write_en(par_done_reg16_write_en),
      .clk(clk),
      .out(par_done_reg16_out),
      .done(par_done_reg16_done)
  );
  
  std_reg #(1) par_reset4 (
      .in(par_reset4_in),
      .write_en(par_reset4_write_en),
      .clk(clk),
      .out(par_reset4_out),
      .done(par_reset4_done)
  );
  
  std_reg #(1) par_done_reg17 (
      .in(par_done_reg17_in),
      .write_en(par_done_reg17_write_en),
      .clk(clk),
      .out(par_done_reg17_out),
      .done(par_done_reg17_done)
  );
  
  std_reg #(1) par_done_reg18 (
      .in(par_done_reg18_in),
      .write_en(par_done_reg18_write_en),
      .clk(clk),
      .out(par_done_reg18_out),
      .done(par_done_reg18_done)
  );
  
  std_reg #(1) par_done_reg19 (
      .in(par_done_reg19_in),
      .write_en(par_done_reg19_write_en),
      .clk(clk),
      .out(par_done_reg19_out),
      .done(par_done_reg19_done)
  );
  
  std_reg #(1) par_done_reg20 (
      .in(par_done_reg20_in),
      .write_en(par_done_reg20_write_en),
      .clk(clk),
      .out(par_done_reg20_out),
      .done(par_done_reg20_done)
  );
  
  std_reg #(1) par_done_reg21 (
      .in(par_done_reg21_in),
      .write_en(par_done_reg21_write_en),
      .clk(clk),
      .out(par_done_reg21_out),
      .done(par_done_reg21_done)
  );
  
  std_reg #(1) par_done_reg22 (
      .in(par_done_reg22_in),
      .write_en(par_done_reg22_write_en),
      .clk(clk),
      .out(par_done_reg22_out),
      .done(par_done_reg22_done)
  );
  
  std_reg #(1) par_reset5 (
      .in(par_reset5_in),
      .write_en(par_reset5_write_en),
      .clk(clk),
      .out(par_reset5_out),
      .done(par_reset5_done)
  );
  
  std_reg #(1) par_done_reg23 (
      .in(par_done_reg23_in),
      .write_en(par_done_reg23_write_en),
      .clk(clk),
      .out(par_done_reg23_out),
      .done(par_done_reg23_done)
  );
  
  std_reg #(1) par_done_reg24 (
      .in(par_done_reg24_in),
      .write_en(par_done_reg24_write_en),
      .clk(clk),
      .out(par_done_reg24_out),
      .done(par_done_reg24_done)
  );
  
  std_reg #(1) par_done_reg25 (
      .in(par_done_reg25_in),
      .write_en(par_done_reg25_write_en),
      .clk(clk),
      .out(par_done_reg25_out),
      .done(par_done_reg25_done)
  );
  
  std_reg #(1) par_done_reg26 (
      .in(par_done_reg26_in),
      .write_en(par_done_reg26_write_en),
      .clk(clk),
      .out(par_done_reg26_out),
      .done(par_done_reg26_done)
  );
  
  std_reg #(1) par_done_reg27 (
      .in(par_done_reg27_in),
      .write_en(par_done_reg27_write_en),
      .clk(clk),
      .out(par_done_reg27_out),
      .done(par_done_reg27_done)
  );
  
  std_reg #(1) par_done_reg28 (
      .in(par_done_reg28_in),
      .write_en(par_done_reg28_write_en),
      .clk(clk),
      .out(par_done_reg28_out),
      .done(par_done_reg28_done)
  );
  
  std_reg #(1) par_done_reg29 (
      .in(par_done_reg29_in),
      .write_en(par_done_reg29_write_en),
      .clk(clk),
      .out(par_done_reg29_out),
      .done(par_done_reg29_done)
  );
  
  std_reg #(1) par_done_reg30 (
      .in(par_done_reg30_in),
      .write_en(par_done_reg30_write_en),
      .clk(clk),
      .out(par_done_reg30_out),
      .done(par_done_reg30_done)
  );
  
  std_reg #(1) par_done_reg31 (
      .in(par_done_reg31_in),
      .write_en(par_done_reg31_write_en),
      .clk(clk),
      .out(par_done_reg31_out),
      .done(par_done_reg31_done)
  );
  
  std_reg #(1) par_reset6 (
      .in(par_reset6_in),
      .write_en(par_reset6_write_en),
      .clk(clk),
      .out(par_reset6_out),
      .done(par_reset6_done)
  );
  
  std_reg #(1) par_done_reg32 (
      .in(par_done_reg32_in),
      .write_en(par_done_reg32_write_en),
      .clk(clk),
      .out(par_done_reg32_out),
      .done(par_done_reg32_done)
  );
  
  std_reg #(1) par_done_reg33 (
      .in(par_done_reg33_in),
      .write_en(par_done_reg33_write_en),
      .clk(clk),
      .out(par_done_reg33_out),
      .done(par_done_reg33_done)
  );
  
  std_reg #(1) par_done_reg34 (
      .in(par_done_reg34_in),
      .write_en(par_done_reg34_write_en),
      .clk(clk),
      .out(par_done_reg34_out),
      .done(par_done_reg34_done)
  );
  
  std_reg #(1) par_done_reg35 (
      .in(par_done_reg35_in),
      .write_en(par_done_reg35_write_en),
      .clk(clk),
      .out(par_done_reg35_out),
      .done(par_done_reg35_done)
  );
  
  std_reg #(1) par_done_reg36 (
      .in(par_done_reg36_in),
      .write_en(par_done_reg36_write_en),
      .clk(clk),
      .out(par_done_reg36_out),
      .done(par_done_reg36_done)
  );
  
  std_reg #(1) par_done_reg37 (
      .in(par_done_reg37_in),
      .write_en(par_done_reg37_write_en),
      .clk(clk),
      .out(par_done_reg37_out),
      .done(par_done_reg37_done)
  );
  
  std_reg #(1) par_done_reg38 (
      .in(par_done_reg38_in),
      .write_en(par_done_reg38_write_en),
      .clk(clk),
      .out(par_done_reg38_out),
      .done(par_done_reg38_done)
  );
  
  std_reg #(1) par_done_reg39 (
      .in(par_done_reg39_in),
      .write_en(par_done_reg39_write_en),
      .clk(clk),
      .out(par_done_reg39_out),
      .done(par_done_reg39_done)
  );
  
  std_reg #(1) par_done_reg40 (
      .in(par_done_reg40_in),
      .write_en(par_done_reg40_write_en),
      .clk(clk),
      .out(par_done_reg40_out),
      .done(par_done_reg40_done)
  );
  
  std_reg #(1) par_done_reg41 (
      .in(par_done_reg41_in),
      .write_en(par_done_reg41_write_en),
      .clk(clk),
      .out(par_done_reg41_out),
      .done(par_done_reg41_done)
  );
  
  std_reg #(1) par_done_reg42 (
      .in(par_done_reg42_in),
      .write_en(par_done_reg42_write_en),
      .clk(clk),
      .out(par_done_reg42_out),
      .done(par_done_reg42_done)
  );
  
  std_reg #(1) par_done_reg43 (
      .in(par_done_reg43_in),
      .write_en(par_done_reg43_write_en),
      .clk(clk),
      .out(par_done_reg43_out),
      .done(par_done_reg43_done)
  );
  
  std_reg #(1) par_reset7 (
      .in(par_reset7_in),
      .write_en(par_reset7_write_en),
      .clk(clk),
      .out(par_reset7_out),
      .done(par_reset7_done)
  );
  
  std_reg #(1) par_done_reg44 (
      .in(par_done_reg44_in),
      .write_en(par_done_reg44_write_en),
      .clk(clk),
      .out(par_done_reg44_out),
      .done(par_done_reg44_done)
  );
  
  std_reg #(1) par_done_reg45 (
      .in(par_done_reg45_in),
      .write_en(par_done_reg45_write_en),
      .clk(clk),
      .out(par_done_reg45_out),
      .done(par_done_reg45_done)
  );
  
  std_reg #(1) par_done_reg46 (
      .in(par_done_reg46_in),
      .write_en(par_done_reg46_write_en),
      .clk(clk),
      .out(par_done_reg46_out),
      .done(par_done_reg46_done)
  );
  
  std_reg #(1) par_done_reg47 (
      .in(par_done_reg47_in),
      .write_en(par_done_reg47_write_en),
      .clk(clk),
      .out(par_done_reg47_out),
      .done(par_done_reg47_done)
  );
  
  std_reg #(1) par_done_reg48 (
      .in(par_done_reg48_in),
      .write_en(par_done_reg48_write_en),
      .clk(clk),
      .out(par_done_reg48_out),
      .done(par_done_reg48_done)
  );
  
  std_reg #(1) par_done_reg49 (
      .in(par_done_reg49_in),
      .write_en(par_done_reg49_write_en),
      .clk(clk),
      .out(par_done_reg49_out),
      .done(par_done_reg49_done)
  );
  
  std_reg #(1) par_done_reg50 (
      .in(par_done_reg50_in),
      .write_en(par_done_reg50_write_en),
      .clk(clk),
      .out(par_done_reg50_out),
      .done(par_done_reg50_done)
  );
  
  std_reg #(1) par_done_reg51 (
      .in(par_done_reg51_in),
      .write_en(par_done_reg51_write_en),
      .clk(clk),
      .out(par_done_reg51_out),
      .done(par_done_reg51_done)
  );
  
  std_reg #(1) par_done_reg52 (
      .in(par_done_reg52_in),
      .write_en(par_done_reg52_write_en),
      .clk(clk),
      .out(par_done_reg52_out),
      .done(par_done_reg52_done)
  );
  
  std_reg #(1) par_done_reg53 (
      .in(par_done_reg53_in),
      .write_en(par_done_reg53_write_en),
      .clk(clk),
      .out(par_done_reg53_out),
      .done(par_done_reg53_done)
  );
  
  std_reg #(1) par_done_reg54 (
      .in(par_done_reg54_in),
      .write_en(par_done_reg54_write_en),
      .clk(clk),
      .out(par_done_reg54_out),
      .done(par_done_reg54_done)
  );
  
  std_reg #(1) par_done_reg55 (
      .in(par_done_reg55_in),
      .write_en(par_done_reg55_write_en),
      .clk(clk),
      .out(par_done_reg55_out),
      .done(par_done_reg55_done)
  );
  
  std_reg #(1) par_done_reg56 (
      .in(par_done_reg56_in),
      .write_en(par_done_reg56_write_en),
      .clk(clk),
      .out(par_done_reg56_out),
      .done(par_done_reg56_done)
  );
  
  std_reg #(1) par_done_reg57 (
      .in(par_done_reg57_in),
      .write_en(par_done_reg57_write_en),
      .clk(clk),
      .out(par_done_reg57_out),
      .done(par_done_reg57_done)
  );
  
  std_reg #(1) par_reset8 (
      .in(par_reset8_in),
      .write_en(par_reset8_write_en),
      .clk(clk),
      .out(par_reset8_out),
      .done(par_reset8_done)
  );
  
  std_reg #(1) par_done_reg58 (
      .in(par_done_reg58_in),
      .write_en(par_done_reg58_write_en),
      .clk(clk),
      .out(par_done_reg58_out),
      .done(par_done_reg58_done)
  );
  
  std_reg #(1) par_done_reg59 (
      .in(par_done_reg59_in),
      .write_en(par_done_reg59_write_en),
      .clk(clk),
      .out(par_done_reg59_out),
      .done(par_done_reg59_done)
  );
  
  std_reg #(1) par_done_reg60 (
      .in(par_done_reg60_in),
      .write_en(par_done_reg60_write_en),
      .clk(clk),
      .out(par_done_reg60_out),
      .done(par_done_reg60_done)
  );
  
  std_reg #(1) par_done_reg61 (
      .in(par_done_reg61_in),
      .write_en(par_done_reg61_write_en),
      .clk(clk),
      .out(par_done_reg61_out),
      .done(par_done_reg61_done)
  );
  
  std_reg #(1) par_done_reg62 (
      .in(par_done_reg62_in),
      .write_en(par_done_reg62_write_en),
      .clk(clk),
      .out(par_done_reg62_out),
      .done(par_done_reg62_done)
  );
  
  std_reg #(1) par_done_reg63 (
      .in(par_done_reg63_in),
      .write_en(par_done_reg63_write_en),
      .clk(clk),
      .out(par_done_reg63_out),
      .done(par_done_reg63_done)
  );
  
  std_reg #(1) par_done_reg64 (
      .in(par_done_reg64_in),
      .write_en(par_done_reg64_write_en),
      .clk(clk),
      .out(par_done_reg64_out),
      .done(par_done_reg64_done)
  );
  
  std_reg #(1) par_done_reg65 (
      .in(par_done_reg65_in),
      .write_en(par_done_reg65_write_en),
      .clk(clk),
      .out(par_done_reg65_out),
      .done(par_done_reg65_done)
  );
  
  std_reg #(1) par_done_reg66 (
      .in(par_done_reg66_in),
      .write_en(par_done_reg66_write_en),
      .clk(clk),
      .out(par_done_reg66_out),
      .done(par_done_reg66_done)
  );
  
  std_reg #(1) par_done_reg67 (
      .in(par_done_reg67_in),
      .write_en(par_done_reg67_write_en),
      .clk(clk),
      .out(par_done_reg67_out),
      .done(par_done_reg67_done)
  );
  
  std_reg #(1) par_done_reg68 (
      .in(par_done_reg68_in),
      .write_en(par_done_reg68_write_en),
      .clk(clk),
      .out(par_done_reg68_out),
      .done(par_done_reg68_done)
  );
  
  std_reg #(1) par_done_reg69 (
      .in(par_done_reg69_in),
      .write_en(par_done_reg69_write_en),
      .clk(clk),
      .out(par_done_reg69_out),
      .done(par_done_reg69_done)
  );
  
  std_reg #(1) par_done_reg70 (
      .in(par_done_reg70_in),
      .write_en(par_done_reg70_write_en),
      .clk(clk),
      .out(par_done_reg70_out),
      .done(par_done_reg70_done)
  );
  
  std_reg #(1) par_done_reg71 (
      .in(par_done_reg71_in),
      .write_en(par_done_reg71_write_en),
      .clk(clk),
      .out(par_done_reg71_out),
      .done(par_done_reg71_done)
  );
  
  std_reg #(1) par_done_reg72 (
      .in(par_done_reg72_in),
      .write_en(par_done_reg72_write_en),
      .clk(clk),
      .out(par_done_reg72_out),
      .done(par_done_reg72_done)
  );
  
  std_reg #(1) par_done_reg73 (
      .in(par_done_reg73_in),
      .write_en(par_done_reg73_write_en),
      .clk(clk),
      .out(par_done_reg73_out),
      .done(par_done_reg73_done)
  );
  
  std_reg #(1) par_done_reg74 (
      .in(par_done_reg74_in),
      .write_en(par_done_reg74_write_en),
      .clk(clk),
      .out(par_done_reg74_out),
      .done(par_done_reg74_done)
  );
  
  std_reg #(1) par_done_reg75 (
      .in(par_done_reg75_in),
      .write_en(par_done_reg75_write_en),
      .clk(clk),
      .out(par_done_reg75_out),
      .done(par_done_reg75_done)
  );
  
  std_reg #(1) par_done_reg76 (
      .in(par_done_reg76_in),
      .write_en(par_done_reg76_write_en),
      .clk(clk),
      .out(par_done_reg76_out),
      .done(par_done_reg76_done)
  );
  
  std_reg #(1) par_done_reg77 (
      .in(par_done_reg77_in),
      .write_en(par_done_reg77_write_en),
      .clk(clk),
      .out(par_done_reg77_out),
      .done(par_done_reg77_done)
  );
  
  std_reg #(1) par_reset9 (
      .in(par_reset9_in),
      .write_en(par_reset9_write_en),
      .clk(clk),
      .out(par_reset9_out),
      .done(par_reset9_done)
  );
  
  std_reg #(1) par_done_reg78 (
      .in(par_done_reg78_in),
      .write_en(par_done_reg78_write_en),
      .clk(clk),
      .out(par_done_reg78_out),
      .done(par_done_reg78_done)
  );
  
  std_reg #(1) par_done_reg79 (
      .in(par_done_reg79_in),
      .write_en(par_done_reg79_write_en),
      .clk(clk),
      .out(par_done_reg79_out),
      .done(par_done_reg79_done)
  );
  
  std_reg #(1) par_done_reg80 (
      .in(par_done_reg80_in),
      .write_en(par_done_reg80_write_en),
      .clk(clk),
      .out(par_done_reg80_out),
      .done(par_done_reg80_done)
  );
  
  std_reg #(1) par_done_reg81 (
      .in(par_done_reg81_in),
      .write_en(par_done_reg81_write_en),
      .clk(clk),
      .out(par_done_reg81_out),
      .done(par_done_reg81_done)
  );
  
  std_reg #(1) par_done_reg82 (
      .in(par_done_reg82_in),
      .write_en(par_done_reg82_write_en),
      .clk(clk),
      .out(par_done_reg82_out),
      .done(par_done_reg82_done)
  );
  
  std_reg #(1) par_done_reg83 (
      .in(par_done_reg83_in),
      .write_en(par_done_reg83_write_en),
      .clk(clk),
      .out(par_done_reg83_out),
      .done(par_done_reg83_done)
  );
  
  std_reg #(1) par_done_reg84 (
      .in(par_done_reg84_in),
      .write_en(par_done_reg84_write_en),
      .clk(clk),
      .out(par_done_reg84_out),
      .done(par_done_reg84_done)
  );
  
  std_reg #(1) par_done_reg85 (
      .in(par_done_reg85_in),
      .write_en(par_done_reg85_write_en),
      .clk(clk),
      .out(par_done_reg85_out),
      .done(par_done_reg85_done)
  );
  
  std_reg #(1) par_done_reg86 (
      .in(par_done_reg86_in),
      .write_en(par_done_reg86_write_en),
      .clk(clk),
      .out(par_done_reg86_out),
      .done(par_done_reg86_done)
  );
  
  std_reg #(1) par_done_reg87 (
      .in(par_done_reg87_in),
      .write_en(par_done_reg87_write_en),
      .clk(clk),
      .out(par_done_reg87_out),
      .done(par_done_reg87_done)
  );
  
  std_reg #(1) par_done_reg88 (
      .in(par_done_reg88_in),
      .write_en(par_done_reg88_write_en),
      .clk(clk),
      .out(par_done_reg88_out),
      .done(par_done_reg88_done)
  );
  
  std_reg #(1) par_done_reg89 (
      .in(par_done_reg89_in),
      .write_en(par_done_reg89_write_en),
      .clk(clk),
      .out(par_done_reg89_out),
      .done(par_done_reg89_done)
  );
  
  std_reg #(1) par_done_reg90 (
      .in(par_done_reg90_in),
      .write_en(par_done_reg90_write_en),
      .clk(clk),
      .out(par_done_reg90_out),
      .done(par_done_reg90_done)
  );
  
  std_reg #(1) par_done_reg91 (
      .in(par_done_reg91_in),
      .write_en(par_done_reg91_write_en),
      .clk(clk),
      .out(par_done_reg91_out),
      .done(par_done_reg91_done)
  );
  
  std_reg #(1) par_done_reg92 (
      .in(par_done_reg92_in),
      .write_en(par_done_reg92_write_en),
      .clk(clk),
      .out(par_done_reg92_out),
      .done(par_done_reg92_done)
  );
  
  std_reg #(1) par_done_reg93 (
      .in(par_done_reg93_in),
      .write_en(par_done_reg93_write_en),
      .clk(clk),
      .out(par_done_reg93_out),
      .done(par_done_reg93_done)
  );
  
  std_reg #(1) par_reset10 (
      .in(par_reset10_in),
      .write_en(par_reset10_write_en),
      .clk(clk),
      .out(par_reset10_out),
      .done(par_reset10_done)
  );
  
  std_reg #(1) par_done_reg94 (
      .in(par_done_reg94_in),
      .write_en(par_done_reg94_write_en),
      .clk(clk),
      .out(par_done_reg94_out),
      .done(par_done_reg94_done)
  );
  
  std_reg #(1) par_done_reg95 (
      .in(par_done_reg95_in),
      .write_en(par_done_reg95_write_en),
      .clk(clk),
      .out(par_done_reg95_out),
      .done(par_done_reg95_done)
  );
  
  std_reg #(1) par_done_reg96 (
      .in(par_done_reg96_in),
      .write_en(par_done_reg96_write_en),
      .clk(clk),
      .out(par_done_reg96_out),
      .done(par_done_reg96_done)
  );
  
  std_reg #(1) par_done_reg97 (
      .in(par_done_reg97_in),
      .write_en(par_done_reg97_write_en),
      .clk(clk),
      .out(par_done_reg97_out),
      .done(par_done_reg97_done)
  );
  
  std_reg #(1) par_done_reg98 (
      .in(par_done_reg98_in),
      .write_en(par_done_reg98_write_en),
      .clk(clk),
      .out(par_done_reg98_out),
      .done(par_done_reg98_done)
  );
  
  std_reg #(1) par_done_reg99 (
      .in(par_done_reg99_in),
      .write_en(par_done_reg99_write_en),
      .clk(clk),
      .out(par_done_reg99_out),
      .done(par_done_reg99_done)
  );
  
  std_reg #(1) par_done_reg100 (
      .in(par_done_reg100_in),
      .write_en(par_done_reg100_write_en),
      .clk(clk),
      .out(par_done_reg100_out),
      .done(par_done_reg100_done)
  );
  
  std_reg #(1) par_done_reg101 (
      .in(par_done_reg101_in),
      .write_en(par_done_reg101_write_en),
      .clk(clk),
      .out(par_done_reg101_out),
      .done(par_done_reg101_done)
  );
  
  std_reg #(1) par_done_reg102 (
      .in(par_done_reg102_in),
      .write_en(par_done_reg102_write_en),
      .clk(clk),
      .out(par_done_reg102_out),
      .done(par_done_reg102_done)
  );
  
  std_reg #(1) par_done_reg103 (
      .in(par_done_reg103_in),
      .write_en(par_done_reg103_write_en),
      .clk(clk),
      .out(par_done_reg103_out),
      .done(par_done_reg103_done)
  );
  
  std_reg #(1) par_done_reg104 (
      .in(par_done_reg104_in),
      .write_en(par_done_reg104_write_en),
      .clk(clk),
      .out(par_done_reg104_out),
      .done(par_done_reg104_done)
  );
  
  std_reg #(1) par_done_reg105 (
      .in(par_done_reg105_in),
      .write_en(par_done_reg105_write_en),
      .clk(clk),
      .out(par_done_reg105_out),
      .done(par_done_reg105_done)
  );
  
  std_reg #(1) par_done_reg106 (
      .in(par_done_reg106_in),
      .write_en(par_done_reg106_write_en),
      .clk(clk),
      .out(par_done_reg106_out),
      .done(par_done_reg106_done)
  );
  
  std_reg #(1) par_done_reg107 (
      .in(par_done_reg107_in),
      .write_en(par_done_reg107_write_en),
      .clk(clk),
      .out(par_done_reg107_out),
      .done(par_done_reg107_done)
  );
  
  std_reg #(1) par_done_reg108 (
      .in(par_done_reg108_in),
      .write_en(par_done_reg108_write_en),
      .clk(clk),
      .out(par_done_reg108_out),
      .done(par_done_reg108_done)
  );
  
  std_reg #(1) par_done_reg109 (
      .in(par_done_reg109_in),
      .write_en(par_done_reg109_write_en),
      .clk(clk),
      .out(par_done_reg109_out),
      .done(par_done_reg109_done)
  );
  
  std_reg #(1) par_done_reg110 (
      .in(par_done_reg110_in),
      .write_en(par_done_reg110_write_en),
      .clk(clk),
      .out(par_done_reg110_out),
      .done(par_done_reg110_done)
  );
  
  std_reg #(1) par_done_reg111 (
      .in(par_done_reg111_in),
      .write_en(par_done_reg111_write_en),
      .clk(clk),
      .out(par_done_reg111_out),
      .done(par_done_reg111_done)
  );
  
  std_reg #(1) par_done_reg112 (
      .in(par_done_reg112_in),
      .write_en(par_done_reg112_write_en),
      .clk(clk),
      .out(par_done_reg112_out),
      .done(par_done_reg112_done)
  );
  
  std_reg #(1) par_done_reg113 (
      .in(par_done_reg113_in),
      .write_en(par_done_reg113_write_en),
      .clk(clk),
      .out(par_done_reg113_out),
      .done(par_done_reg113_done)
  );
  
  std_reg #(1) par_done_reg114 (
      .in(par_done_reg114_in),
      .write_en(par_done_reg114_write_en),
      .clk(clk),
      .out(par_done_reg114_out),
      .done(par_done_reg114_done)
  );
  
  std_reg #(1) par_done_reg115 (
      .in(par_done_reg115_in),
      .write_en(par_done_reg115_write_en),
      .clk(clk),
      .out(par_done_reg115_out),
      .done(par_done_reg115_done)
  );
  
  std_reg #(1) par_done_reg116 (
      .in(par_done_reg116_in),
      .write_en(par_done_reg116_write_en),
      .clk(clk),
      .out(par_done_reg116_out),
      .done(par_done_reg116_done)
  );
  
  std_reg #(1) par_done_reg117 (
      .in(par_done_reg117_in),
      .write_en(par_done_reg117_write_en),
      .clk(clk),
      .out(par_done_reg117_out),
      .done(par_done_reg117_done)
  );
  
  std_reg #(1) par_reset11 (
      .in(par_reset11_in),
      .write_en(par_reset11_write_en),
      .clk(clk),
      .out(par_reset11_out),
      .done(par_reset11_done)
  );
  
  std_reg #(1) par_done_reg118 (
      .in(par_done_reg118_in),
      .write_en(par_done_reg118_write_en),
      .clk(clk),
      .out(par_done_reg118_out),
      .done(par_done_reg118_done)
  );
  
  std_reg #(1) par_done_reg119 (
      .in(par_done_reg119_in),
      .write_en(par_done_reg119_write_en),
      .clk(clk),
      .out(par_done_reg119_out),
      .done(par_done_reg119_done)
  );
  
  std_reg #(1) par_done_reg120 (
      .in(par_done_reg120_in),
      .write_en(par_done_reg120_write_en),
      .clk(clk),
      .out(par_done_reg120_out),
      .done(par_done_reg120_done)
  );
  
  std_reg #(1) par_done_reg121 (
      .in(par_done_reg121_in),
      .write_en(par_done_reg121_write_en),
      .clk(clk),
      .out(par_done_reg121_out),
      .done(par_done_reg121_done)
  );
  
  std_reg #(1) par_done_reg122 (
      .in(par_done_reg122_in),
      .write_en(par_done_reg122_write_en),
      .clk(clk),
      .out(par_done_reg122_out),
      .done(par_done_reg122_done)
  );
  
  std_reg #(1) par_done_reg123 (
      .in(par_done_reg123_in),
      .write_en(par_done_reg123_write_en),
      .clk(clk),
      .out(par_done_reg123_out),
      .done(par_done_reg123_done)
  );
  
  std_reg #(1) par_done_reg124 (
      .in(par_done_reg124_in),
      .write_en(par_done_reg124_write_en),
      .clk(clk),
      .out(par_done_reg124_out),
      .done(par_done_reg124_done)
  );
  
  std_reg #(1) par_done_reg125 (
      .in(par_done_reg125_in),
      .write_en(par_done_reg125_write_en),
      .clk(clk),
      .out(par_done_reg125_out),
      .done(par_done_reg125_done)
  );
  
  std_reg #(1) par_done_reg126 (
      .in(par_done_reg126_in),
      .write_en(par_done_reg126_write_en),
      .clk(clk),
      .out(par_done_reg126_out),
      .done(par_done_reg126_done)
  );
  
  std_reg #(1) par_done_reg127 (
      .in(par_done_reg127_in),
      .write_en(par_done_reg127_write_en),
      .clk(clk),
      .out(par_done_reg127_out),
      .done(par_done_reg127_done)
  );
  
  std_reg #(1) par_done_reg128 (
      .in(par_done_reg128_in),
      .write_en(par_done_reg128_write_en),
      .clk(clk),
      .out(par_done_reg128_out),
      .done(par_done_reg128_done)
  );
  
  std_reg #(1) par_done_reg129 (
      .in(par_done_reg129_in),
      .write_en(par_done_reg129_write_en),
      .clk(clk),
      .out(par_done_reg129_out),
      .done(par_done_reg129_done)
  );
  
  std_reg #(1) par_done_reg130 (
      .in(par_done_reg130_in),
      .write_en(par_done_reg130_write_en),
      .clk(clk),
      .out(par_done_reg130_out),
      .done(par_done_reg130_done)
  );
  
  std_reg #(1) par_done_reg131 (
      .in(par_done_reg131_in),
      .write_en(par_done_reg131_write_en),
      .clk(clk),
      .out(par_done_reg131_out),
      .done(par_done_reg131_done)
  );
  
  std_reg #(1) par_done_reg132 (
      .in(par_done_reg132_in),
      .write_en(par_done_reg132_write_en),
      .clk(clk),
      .out(par_done_reg132_out),
      .done(par_done_reg132_done)
  );
  
  std_reg #(1) par_done_reg133 (
      .in(par_done_reg133_in),
      .write_en(par_done_reg133_write_en),
      .clk(clk),
      .out(par_done_reg133_out),
      .done(par_done_reg133_done)
  );
  
  std_reg #(1) par_reset12 (
      .in(par_reset12_in),
      .write_en(par_reset12_write_en),
      .clk(clk),
      .out(par_reset12_out),
      .done(par_reset12_done)
  );
  
  std_reg #(1) par_done_reg134 (
      .in(par_done_reg134_in),
      .write_en(par_done_reg134_write_en),
      .clk(clk),
      .out(par_done_reg134_out),
      .done(par_done_reg134_done)
  );
  
  std_reg #(1) par_done_reg135 (
      .in(par_done_reg135_in),
      .write_en(par_done_reg135_write_en),
      .clk(clk),
      .out(par_done_reg135_out),
      .done(par_done_reg135_done)
  );
  
  std_reg #(1) par_done_reg136 (
      .in(par_done_reg136_in),
      .write_en(par_done_reg136_write_en),
      .clk(clk),
      .out(par_done_reg136_out),
      .done(par_done_reg136_done)
  );
  
  std_reg #(1) par_done_reg137 (
      .in(par_done_reg137_in),
      .write_en(par_done_reg137_write_en),
      .clk(clk),
      .out(par_done_reg137_out),
      .done(par_done_reg137_done)
  );
  
  std_reg #(1) par_done_reg138 (
      .in(par_done_reg138_in),
      .write_en(par_done_reg138_write_en),
      .clk(clk),
      .out(par_done_reg138_out),
      .done(par_done_reg138_done)
  );
  
  std_reg #(1) par_done_reg139 (
      .in(par_done_reg139_in),
      .write_en(par_done_reg139_write_en),
      .clk(clk),
      .out(par_done_reg139_out),
      .done(par_done_reg139_done)
  );
  
  std_reg #(1) par_done_reg140 (
      .in(par_done_reg140_in),
      .write_en(par_done_reg140_write_en),
      .clk(clk),
      .out(par_done_reg140_out),
      .done(par_done_reg140_done)
  );
  
  std_reg #(1) par_done_reg141 (
      .in(par_done_reg141_in),
      .write_en(par_done_reg141_write_en),
      .clk(clk),
      .out(par_done_reg141_out),
      .done(par_done_reg141_done)
  );
  
  std_reg #(1) par_done_reg142 (
      .in(par_done_reg142_in),
      .write_en(par_done_reg142_write_en),
      .clk(clk),
      .out(par_done_reg142_out),
      .done(par_done_reg142_done)
  );
  
  std_reg #(1) par_done_reg143 (
      .in(par_done_reg143_in),
      .write_en(par_done_reg143_write_en),
      .clk(clk),
      .out(par_done_reg143_out),
      .done(par_done_reg143_done)
  );
  
  std_reg #(1) par_done_reg144 (
      .in(par_done_reg144_in),
      .write_en(par_done_reg144_write_en),
      .clk(clk),
      .out(par_done_reg144_out),
      .done(par_done_reg144_done)
  );
  
  std_reg #(1) par_done_reg145 (
      .in(par_done_reg145_in),
      .write_en(par_done_reg145_write_en),
      .clk(clk),
      .out(par_done_reg145_out),
      .done(par_done_reg145_done)
  );
  
  std_reg #(1) par_done_reg146 (
      .in(par_done_reg146_in),
      .write_en(par_done_reg146_write_en),
      .clk(clk),
      .out(par_done_reg146_out),
      .done(par_done_reg146_done)
  );
  
  std_reg #(1) par_done_reg147 (
      .in(par_done_reg147_in),
      .write_en(par_done_reg147_write_en),
      .clk(clk),
      .out(par_done_reg147_out),
      .done(par_done_reg147_done)
  );
  
  std_reg #(1) par_done_reg148 (
      .in(par_done_reg148_in),
      .write_en(par_done_reg148_write_en),
      .clk(clk),
      .out(par_done_reg148_out),
      .done(par_done_reg148_done)
  );
  
  std_reg #(1) par_done_reg149 (
      .in(par_done_reg149_in),
      .write_en(par_done_reg149_write_en),
      .clk(clk),
      .out(par_done_reg149_out),
      .done(par_done_reg149_done)
  );
  
  std_reg #(1) par_done_reg150 (
      .in(par_done_reg150_in),
      .write_en(par_done_reg150_write_en),
      .clk(clk),
      .out(par_done_reg150_out),
      .done(par_done_reg150_done)
  );
  
  std_reg #(1) par_done_reg151 (
      .in(par_done_reg151_in),
      .write_en(par_done_reg151_write_en),
      .clk(clk),
      .out(par_done_reg151_out),
      .done(par_done_reg151_done)
  );
  
  std_reg #(1) par_done_reg152 (
      .in(par_done_reg152_in),
      .write_en(par_done_reg152_write_en),
      .clk(clk),
      .out(par_done_reg152_out),
      .done(par_done_reg152_done)
  );
  
  std_reg #(1) par_done_reg153 (
      .in(par_done_reg153_in),
      .write_en(par_done_reg153_write_en),
      .clk(clk),
      .out(par_done_reg153_out),
      .done(par_done_reg153_done)
  );
  
  std_reg #(1) par_done_reg154 (
      .in(par_done_reg154_in),
      .write_en(par_done_reg154_write_en),
      .clk(clk),
      .out(par_done_reg154_out),
      .done(par_done_reg154_done)
  );
  
  std_reg #(1) par_done_reg155 (
      .in(par_done_reg155_in),
      .write_en(par_done_reg155_write_en),
      .clk(clk),
      .out(par_done_reg155_out),
      .done(par_done_reg155_done)
  );
  
  std_reg #(1) par_done_reg156 (
      .in(par_done_reg156_in),
      .write_en(par_done_reg156_write_en),
      .clk(clk),
      .out(par_done_reg156_out),
      .done(par_done_reg156_done)
  );
  
  std_reg #(1) par_done_reg157 (
      .in(par_done_reg157_in),
      .write_en(par_done_reg157_write_en),
      .clk(clk),
      .out(par_done_reg157_out),
      .done(par_done_reg157_done)
  );
  
  std_reg #(1) par_reset13 (
      .in(par_reset13_in),
      .write_en(par_reset13_write_en),
      .clk(clk),
      .out(par_reset13_out),
      .done(par_reset13_done)
  );
  
  std_reg #(1) par_done_reg158 (
      .in(par_done_reg158_in),
      .write_en(par_done_reg158_write_en),
      .clk(clk),
      .out(par_done_reg158_out),
      .done(par_done_reg158_done)
  );
  
  std_reg #(1) par_done_reg159 (
      .in(par_done_reg159_in),
      .write_en(par_done_reg159_write_en),
      .clk(clk),
      .out(par_done_reg159_out),
      .done(par_done_reg159_done)
  );
  
  std_reg #(1) par_done_reg160 (
      .in(par_done_reg160_in),
      .write_en(par_done_reg160_write_en),
      .clk(clk),
      .out(par_done_reg160_out),
      .done(par_done_reg160_done)
  );
  
  std_reg #(1) par_done_reg161 (
      .in(par_done_reg161_in),
      .write_en(par_done_reg161_write_en),
      .clk(clk),
      .out(par_done_reg161_out),
      .done(par_done_reg161_done)
  );
  
  std_reg #(1) par_done_reg162 (
      .in(par_done_reg162_in),
      .write_en(par_done_reg162_write_en),
      .clk(clk),
      .out(par_done_reg162_out),
      .done(par_done_reg162_done)
  );
  
  std_reg #(1) par_done_reg163 (
      .in(par_done_reg163_in),
      .write_en(par_done_reg163_write_en),
      .clk(clk),
      .out(par_done_reg163_out),
      .done(par_done_reg163_done)
  );
  
  std_reg #(1) par_done_reg164 (
      .in(par_done_reg164_in),
      .write_en(par_done_reg164_write_en),
      .clk(clk),
      .out(par_done_reg164_out),
      .done(par_done_reg164_done)
  );
  
  std_reg #(1) par_done_reg165 (
      .in(par_done_reg165_in),
      .write_en(par_done_reg165_write_en),
      .clk(clk),
      .out(par_done_reg165_out),
      .done(par_done_reg165_done)
  );
  
  std_reg #(1) par_done_reg166 (
      .in(par_done_reg166_in),
      .write_en(par_done_reg166_write_en),
      .clk(clk),
      .out(par_done_reg166_out),
      .done(par_done_reg166_done)
  );
  
  std_reg #(1) par_done_reg167 (
      .in(par_done_reg167_in),
      .write_en(par_done_reg167_write_en),
      .clk(clk),
      .out(par_done_reg167_out),
      .done(par_done_reg167_done)
  );
  
  std_reg #(1) par_done_reg168 (
      .in(par_done_reg168_in),
      .write_en(par_done_reg168_write_en),
      .clk(clk),
      .out(par_done_reg168_out),
      .done(par_done_reg168_done)
  );
  
  std_reg #(1) par_done_reg169 (
      .in(par_done_reg169_in),
      .write_en(par_done_reg169_write_en),
      .clk(clk),
      .out(par_done_reg169_out),
      .done(par_done_reg169_done)
  );
  
  std_reg #(1) par_done_reg170 (
      .in(par_done_reg170_in),
      .write_en(par_done_reg170_write_en),
      .clk(clk),
      .out(par_done_reg170_out),
      .done(par_done_reg170_done)
  );
  
  std_reg #(1) par_done_reg171 (
      .in(par_done_reg171_in),
      .write_en(par_done_reg171_write_en),
      .clk(clk),
      .out(par_done_reg171_out),
      .done(par_done_reg171_done)
  );
  
  std_reg #(1) par_reset14 (
      .in(par_reset14_in),
      .write_en(par_reset14_write_en),
      .clk(clk),
      .out(par_reset14_out),
      .done(par_reset14_done)
  );
  
  std_reg #(1) par_done_reg172 (
      .in(par_done_reg172_in),
      .write_en(par_done_reg172_write_en),
      .clk(clk),
      .out(par_done_reg172_out),
      .done(par_done_reg172_done)
  );
  
  std_reg #(1) par_done_reg173 (
      .in(par_done_reg173_in),
      .write_en(par_done_reg173_write_en),
      .clk(clk),
      .out(par_done_reg173_out),
      .done(par_done_reg173_done)
  );
  
  std_reg #(1) par_done_reg174 (
      .in(par_done_reg174_in),
      .write_en(par_done_reg174_write_en),
      .clk(clk),
      .out(par_done_reg174_out),
      .done(par_done_reg174_done)
  );
  
  std_reg #(1) par_done_reg175 (
      .in(par_done_reg175_in),
      .write_en(par_done_reg175_write_en),
      .clk(clk),
      .out(par_done_reg175_out),
      .done(par_done_reg175_done)
  );
  
  std_reg #(1) par_done_reg176 (
      .in(par_done_reg176_in),
      .write_en(par_done_reg176_write_en),
      .clk(clk),
      .out(par_done_reg176_out),
      .done(par_done_reg176_done)
  );
  
  std_reg #(1) par_done_reg177 (
      .in(par_done_reg177_in),
      .write_en(par_done_reg177_write_en),
      .clk(clk),
      .out(par_done_reg177_out),
      .done(par_done_reg177_done)
  );
  
  std_reg #(1) par_done_reg178 (
      .in(par_done_reg178_in),
      .write_en(par_done_reg178_write_en),
      .clk(clk),
      .out(par_done_reg178_out),
      .done(par_done_reg178_done)
  );
  
  std_reg #(1) par_done_reg179 (
      .in(par_done_reg179_in),
      .write_en(par_done_reg179_write_en),
      .clk(clk),
      .out(par_done_reg179_out),
      .done(par_done_reg179_done)
  );
  
  std_reg #(1) par_done_reg180 (
      .in(par_done_reg180_in),
      .write_en(par_done_reg180_write_en),
      .clk(clk),
      .out(par_done_reg180_out),
      .done(par_done_reg180_done)
  );
  
  std_reg #(1) par_done_reg181 (
      .in(par_done_reg181_in),
      .write_en(par_done_reg181_write_en),
      .clk(clk),
      .out(par_done_reg181_out),
      .done(par_done_reg181_done)
  );
  
  std_reg #(1) par_done_reg182 (
      .in(par_done_reg182_in),
      .write_en(par_done_reg182_write_en),
      .clk(clk),
      .out(par_done_reg182_out),
      .done(par_done_reg182_done)
  );
  
  std_reg #(1) par_done_reg183 (
      .in(par_done_reg183_in),
      .write_en(par_done_reg183_write_en),
      .clk(clk),
      .out(par_done_reg183_out),
      .done(par_done_reg183_done)
  );
  
  std_reg #(1) par_done_reg184 (
      .in(par_done_reg184_in),
      .write_en(par_done_reg184_write_en),
      .clk(clk),
      .out(par_done_reg184_out),
      .done(par_done_reg184_done)
  );
  
  std_reg #(1) par_done_reg185 (
      .in(par_done_reg185_in),
      .write_en(par_done_reg185_write_en),
      .clk(clk),
      .out(par_done_reg185_out),
      .done(par_done_reg185_done)
  );
  
  std_reg #(1) par_done_reg186 (
      .in(par_done_reg186_in),
      .write_en(par_done_reg186_write_en),
      .clk(clk),
      .out(par_done_reg186_out),
      .done(par_done_reg186_done)
  );
  
  std_reg #(1) par_done_reg187 (
      .in(par_done_reg187_in),
      .write_en(par_done_reg187_write_en),
      .clk(clk),
      .out(par_done_reg187_out),
      .done(par_done_reg187_done)
  );
  
  std_reg #(1) par_done_reg188 (
      .in(par_done_reg188_in),
      .write_en(par_done_reg188_write_en),
      .clk(clk),
      .out(par_done_reg188_out),
      .done(par_done_reg188_done)
  );
  
  std_reg #(1) par_done_reg189 (
      .in(par_done_reg189_in),
      .write_en(par_done_reg189_write_en),
      .clk(clk),
      .out(par_done_reg189_out),
      .done(par_done_reg189_done)
  );
  
  std_reg #(1) par_done_reg190 (
      .in(par_done_reg190_in),
      .write_en(par_done_reg190_write_en),
      .clk(clk),
      .out(par_done_reg190_out),
      .done(par_done_reg190_done)
  );
  
  std_reg #(1) par_done_reg191 (
      .in(par_done_reg191_in),
      .write_en(par_done_reg191_write_en),
      .clk(clk),
      .out(par_done_reg191_out),
      .done(par_done_reg191_done)
  );
  
  std_reg #(1) par_reset15 (
      .in(par_reset15_in),
      .write_en(par_reset15_write_en),
      .clk(clk),
      .out(par_reset15_out),
      .done(par_reset15_done)
  );
  
  std_reg #(1) par_done_reg192 (
      .in(par_done_reg192_in),
      .write_en(par_done_reg192_write_en),
      .clk(clk),
      .out(par_done_reg192_out),
      .done(par_done_reg192_done)
  );
  
  std_reg #(1) par_done_reg193 (
      .in(par_done_reg193_in),
      .write_en(par_done_reg193_write_en),
      .clk(clk),
      .out(par_done_reg193_out),
      .done(par_done_reg193_done)
  );
  
  std_reg #(1) par_done_reg194 (
      .in(par_done_reg194_in),
      .write_en(par_done_reg194_write_en),
      .clk(clk),
      .out(par_done_reg194_out),
      .done(par_done_reg194_done)
  );
  
  std_reg #(1) par_done_reg195 (
      .in(par_done_reg195_in),
      .write_en(par_done_reg195_write_en),
      .clk(clk),
      .out(par_done_reg195_out),
      .done(par_done_reg195_done)
  );
  
  std_reg #(1) par_done_reg196 (
      .in(par_done_reg196_in),
      .write_en(par_done_reg196_write_en),
      .clk(clk),
      .out(par_done_reg196_out),
      .done(par_done_reg196_done)
  );
  
  std_reg #(1) par_done_reg197 (
      .in(par_done_reg197_in),
      .write_en(par_done_reg197_write_en),
      .clk(clk),
      .out(par_done_reg197_out),
      .done(par_done_reg197_done)
  );
  
  std_reg #(1) par_done_reg198 (
      .in(par_done_reg198_in),
      .write_en(par_done_reg198_write_en),
      .clk(clk),
      .out(par_done_reg198_out),
      .done(par_done_reg198_done)
  );
  
  std_reg #(1) par_done_reg199 (
      .in(par_done_reg199_in),
      .write_en(par_done_reg199_write_en),
      .clk(clk),
      .out(par_done_reg199_out),
      .done(par_done_reg199_done)
  );
  
  std_reg #(1) par_done_reg200 (
      .in(par_done_reg200_in),
      .write_en(par_done_reg200_write_en),
      .clk(clk),
      .out(par_done_reg200_out),
      .done(par_done_reg200_done)
  );
  
  std_reg #(1) par_done_reg201 (
      .in(par_done_reg201_in),
      .write_en(par_done_reg201_write_en),
      .clk(clk),
      .out(par_done_reg201_out),
      .done(par_done_reg201_done)
  );
  
  std_reg #(1) par_reset16 (
      .in(par_reset16_in),
      .write_en(par_reset16_write_en),
      .clk(clk),
      .out(par_reset16_out),
      .done(par_reset16_done)
  );
  
  std_reg #(1) par_done_reg202 (
      .in(par_done_reg202_in),
      .write_en(par_done_reg202_write_en),
      .clk(clk),
      .out(par_done_reg202_out),
      .done(par_done_reg202_done)
  );
  
  std_reg #(1) par_done_reg203 (
      .in(par_done_reg203_in),
      .write_en(par_done_reg203_write_en),
      .clk(clk),
      .out(par_done_reg203_out),
      .done(par_done_reg203_done)
  );
  
  std_reg #(1) par_done_reg204 (
      .in(par_done_reg204_in),
      .write_en(par_done_reg204_write_en),
      .clk(clk),
      .out(par_done_reg204_out),
      .done(par_done_reg204_done)
  );
  
  std_reg #(1) par_done_reg205 (
      .in(par_done_reg205_in),
      .write_en(par_done_reg205_write_en),
      .clk(clk),
      .out(par_done_reg205_out),
      .done(par_done_reg205_done)
  );
  
  std_reg #(1) par_done_reg206 (
      .in(par_done_reg206_in),
      .write_en(par_done_reg206_write_en),
      .clk(clk),
      .out(par_done_reg206_out),
      .done(par_done_reg206_done)
  );
  
  std_reg #(1) par_done_reg207 (
      .in(par_done_reg207_in),
      .write_en(par_done_reg207_write_en),
      .clk(clk),
      .out(par_done_reg207_out),
      .done(par_done_reg207_done)
  );
  
  std_reg #(1) par_done_reg208 (
      .in(par_done_reg208_in),
      .write_en(par_done_reg208_write_en),
      .clk(clk),
      .out(par_done_reg208_out),
      .done(par_done_reg208_done)
  );
  
  std_reg #(1) par_done_reg209 (
      .in(par_done_reg209_in),
      .write_en(par_done_reg209_write_en),
      .clk(clk),
      .out(par_done_reg209_out),
      .done(par_done_reg209_done)
  );
  
  std_reg #(1) par_done_reg210 (
      .in(par_done_reg210_in),
      .write_en(par_done_reg210_write_en),
      .clk(clk),
      .out(par_done_reg210_out),
      .done(par_done_reg210_done)
  );
  
  std_reg #(1) par_done_reg211 (
      .in(par_done_reg211_in),
      .write_en(par_done_reg211_write_en),
      .clk(clk),
      .out(par_done_reg211_out),
      .done(par_done_reg211_done)
  );
  
  std_reg #(1) par_done_reg212 (
      .in(par_done_reg212_in),
      .write_en(par_done_reg212_write_en),
      .clk(clk),
      .out(par_done_reg212_out),
      .done(par_done_reg212_done)
  );
  
  std_reg #(1) par_done_reg213 (
      .in(par_done_reg213_in),
      .write_en(par_done_reg213_write_en),
      .clk(clk),
      .out(par_done_reg213_out),
      .done(par_done_reg213_done)
  );
  
  std_reg #(1) par_reset17 (
      .in(par_reset17_in),
      .write_en(par_reset17_write_en),
      .clk(clk),
      .out(par_reset17_out),
      .done(par_reset17_done)
  );
  
  std_reg #(1) par_done_reg214 (
      .in(par_done_reg214_in),
      .write_en(par_done_reg214_write_en),
      .clk(clk),
      .out(par_done_reg214_out),
      .done(par_done_reg214_done)
  );
  
  std_reg #(1) par_done_reg215 (
      .in(par_done_reg215_in),
      .write_en(par_done_reg215_write_en),
      .clk(clk),
      .out(par_done_reg215_out),
      .done(par_done_reg215_done)
  );
  
  std_reg #(1) par_done_reg216 (
      .in(par_done_reg216_in),
      .write_en(par_done_reg216_write_en),
      .clk(clk),
      .out(par_done_reg216_out),
      .done(par_done_reg216_done)
  );
  
  std_reg #(1) par_done_reg217 (
      .in(par_done_reg217_in),
      .write_en(par_done_reg217_write_en),
      .clk(clk),
      .out(par_done_reg217_out),
      .done(par_done_reg217_done)
  );
  
  std_reg #(1) par_done_reg218 (
      .in(par_done_reg218_in),
      .write_en(par_done_reg218_write_en),
      .clk(clk),
      .out(par_done_reg218_out),
      .done(par_done_reg218_done)
  );
  
  std_reg #(1) par_done_reg219 (
      .in(par_done_reg219_in),
      .write_en(par_done_reg219_write_en),
      .clk(clk),
      .out(par_done_reg219_out),
      .done(par_done_reg219_done)
  );
  
  std_reg #(1) par_reset18 (
      .in(par_reset18_in),
      .write_en(par_reset18_write_en),
      .clk(clk),
      .out(par_reset18_out),
      .done(par_reset18_done)
  );
  
  std_reg #(1) par_done_reg220 (
      .in(par_done_reg220_in),
      .write_en(par_done_reg220_write_en),
      .clk(clk),
      .out(par_done_reg220_out),
      .done(par_done_reg220_done)
  );
  
  std_reg #(1) par_done_reg221 (
      .in(par_done_reg221_in),
      .write_en(par_done_reg221_write_en),
      .clk(clk),
      .out(par_done_reg221_out),
      .done(par_done_reg221_done)
  );
  
  std_reg #(1) par_done_reg222 (
      .in(par_done_reg222_in),
      .write_en(par_done_reg222_write_en),
      .clk(clk),
      .out(par_done_reg222_out),
      .done(par_done_reg222_done)
  );
  
  std_reg #(1) par_done_reg223 (
      .in(par_done_reg223_in),
      .write_en(par_done_reg223_write_en),
      .clk(clk),
      .out(par_done_reg223_out),
      .done(par_done_reg223_done)
  );
  
  std_reg #(1) par_done_reg224 (
      .in(par_done_reg224_in),
      .write_en(par_done_reg224_write_en),
      .clk(clk),
      .out(par_done_reg224_out),
      .done(par_done_reg224_done)
  );
  
  std_reg #(1) par_done_reg225 (
      .in(par_done_reg225_in),
      .write_en(par_done_reg225_write_en),
      .clk(clk),
      .out(par_done_reg225_out),
      .done(par_done_reg225_done)
  );
  
  std_reg #(1) par_reset19 (
      .in(par_reset19_in),
      .write_en(par_reset19_write_en),
      .clk(clk),
      .out(par_reset19_out),
      .done(par_reset19_done)
  );
  
  std_reg #(1) par_done_reg226 (
      .in(par_done_reg226_in),
      .write_en(par_done_reg226_write_en),
      .clk(clk),
      .out(par_done_reg226_out),
      .done(par_done_reg226_done)
  );
  
  std_reg #(1) par_done_reg227 (
      .in(par_done_reg227_in),
      .write_en(par_done_reg227_write_en),
      .clk(clk),
      .out(par_done_reg227_out),
      .done(par_done_reg227_done)
  );
  
  std_reg #(1) par_done_reg228 (
      .in(par_done_reg228_in),
      .write_en(par_done_reg228_write_en),
      .clk(clk),
      .out(par_done_reg228_out),
      .done(par_done_reg228_done)
  );
  
  std_reg #(1) par_reset20 (
      .in(par_reset20_in),
      .write_en(par_reset20_write_en),
      .clk(clk),
      .out(par_reset20_out),
      .done(par_reset20_done)
  );
  
  std_reg #(1) par_done_reg229 (
      .in(par_done_reg229_in),
      .write_en(par_done_reg229_write_en),
      .clk(clk),
      .out(par_done_reg229_out),
      .done(par_done_reg229_done)
  );
  
  std_reg #(1) par_done_reg230 (
      .in(par_done_reg230_in),
      .write_en(par_done_reg230_write_en),
      .clk(clk),
      .out(par_done_reg230_out),
      .done(par_done_reg230_done)
  );
  
  std_reg #(1) par_reset21 (
      .in(par_reset21_in),
      .write_en(par_reset21_write_en),
      .clk(clk),
      .out(par_reset21_out),
      .done(par_reset21_done)
  );
  
  std_reg #(1) par_done_reg231 (
      .in(par_done_reg231_in),
      .write_en(par_done_reg231_write_en),
      .clk(clk),
      .out(par_done_reg231_out),
      .done(par_done_reg231_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign done = (fsm0_out == 32'd38) ? 1'd1 : '0;
  assign out_mem_addr0 = (fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go) ? 3'd3 : (fsm0_out == 32'd30 & !out_mem_done & go | fsm0_out == 32'd31 & !out_mem_done & go | fsm0_out == 32'd32 & !out_mem_done & go | fsm0_out == 32'd33 & !out_mem_done & go) ? 3'd2 : (fsm0_out == 32'd22 & !out_mem_done & go | fsm0_out == 32'd23 & !out_mem_done & go | fsm0_out == 32'd24 & !out_mem_done & go | fsm0_out == 32'd25 & !out_mem_done & go) ? 3'd0 : (fsm0_out == 32'd26 & !out_mem_done & go | fsm0_out == 32'd27 & !out_mem_done & go | fsm0_out == 32'd28 & !out_mem_done & go | fsm0_out == 32'd29 & !out_mem_done & go) ? 3'd1 : '0;
  assign out_mem_addr1 = (fsm0_out == 32'd25 & !out_mem_done & go | fsm0_out == 32'd29 & !out_mem_done & go | fsm0_out == 32'd33 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go) ? 3'd3 : (fsm0_out == 32'd24 & !out_mem_done & go | fsm0_out == 32'd28 & !out_mem_done & go | fsm0_out == 32'd32 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go) ? 3'd2 : (fsm0_out == 32'd22 & !out_mem_done & go | fsm0_out == 32'd26 & !out_mem_done & go | fsm0_out == 32'd30 & !out_mem_done & go | fsm0_out == 32'd34 & !out_mem_done & go) ? 3'd0 : (fsm0_out == 32'd23 & !out_mem_done & go | fsm0_out == 32'd27 & !out_mem_done & go | fsm0_out == 32'd31 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go) ? 3'd1 : '0;
  assign out_mem_write_data = (fsm0_out == 32'd37 & !out_mem_done & go) ? pe_33_out : (fsm0_out == 32'd36 & !out_mem_done & go) ? pe_32_out : (fsm0_out == 32'd35 & !out_mem_done & go) ? pe_31_out : (fsm0_out == 32'd34 & !out_mem_done & go) ? pe_30_out : (fsm0_out == 32'd33 & !out_mem_done & go) ? pe_23_out : (fsm0_out == 32'd32 & !out_mem_done & go) ? pe_22_out : (fsm0_out == 32'd31 & !out_mem_done & go) ? pe_21_out : (fsm0_out == 32'd30 & !out_mem_done & go) ? pe_20_out : (fsm0_out == 32'd29 & !out_mem_done & go) ? pe_13_out : (fsm0_out == 32'd28 & !out_mem_done & go) ? pe_12_out : (fsm0_out == 32'd27 & !out_mem_done & go) ? pe_11_out : (fsm0_out == 32'd26 & !out_mem_done & go) ? pe_10_out : (fsm0_out == 32'd25 & !out_mem_done & go) ? pe_03_out : (fsm0_out == 32'd24 & !out_mem_done & go) ? pe_02_out : (fsm0_out == 32'd23 & !out_mem_done & go) ? pe_01_out : (fsm0_out == 32'd22 & !out_mem_done & go) ? pe_00_out : '0;
  assign out_mem_write_en = (fsm0_out == 32'd22 & !out_mem_done & go | fsm0_out == 32'd23 & !out_mem_done & go | fsm0_out == 32'd24 & !out_mem_done & go | fsm0_out == 32'd25 & !out_mem_done & go | fsm0_out == 32'd26 & !out_mem_done & go | fsm0_out == 32'd27 & !out_mem_done & go | fsm0_out == 32'd28 & !out_mem_done & go | fsm0_out == 32'd29 & !out_mem_done & go | fsm0_out == 32'd30 & !out_mem_done & go | fsm0_out == 32'd31 & !out_mem_done & go | fsm0_out == 32'd32 & !out_mem_done & go | fsm0_out == 32'd33 & !out_mem_done & go | fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go) ? 1'd1 : '0;
  assign left_33_read_in = (!(par_done_reg191_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg213_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg225_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg230_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_32_write_out : '0;
  assign left_33_read_write_en = (!(par_done_reg191_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg213_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg225_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg230_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_33_read_in = (!(par_done_reg181_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg207_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg222_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg229_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_23_write_out : '0;
  assign top_33_read_write_en = (!(par_done_reg181_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg207_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg222_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg229_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_33_top = (!(par_done_reg201_out | pe_33_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg219_out | pe_33_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg228_out | pe_33_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg231_out | pe_33_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_33_read_out : '0;
  assign pe_33_left = (!(par_done_reg201_out | pe_33_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg219_out | pe_33_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg228_out | pe_33_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg231_out | pe_33_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_33_read_out : '0;
  assign pe_33_go = (!pe_33_done & (!(par_done_reg201_out | pe_33_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg219_out | pe_33_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg228_out | pe_33_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg231_out | pe_33_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_32_write_in = (pe_32_done & (!(par_done_reg171_out | right_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg200_out | right_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg218_out | right_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg227_out | right_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_32_right : '0;
  assign right_32_write_write_en = (pe_32_done & (!(par_done_reg171_out | right_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg200_out | right_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg218_out | right_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg227_out | right_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_32_read_in = (!(par_done_reg157_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg190_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg212_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg224_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_31_write_out : '0;
  assign left_32_read_write_en = (!(par_done_reg157_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg190_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg212_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg224_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_32_read_in = (!(par_done_reg145_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg180_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg206_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg221_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_22_write_out : '0;
  assign top_32_read_write_en = (!(par_done_reg145_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg180_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg206_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg221_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_32_top = (!(par_done_reg171_out | right_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg200_out | right_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg218_out | right_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg227_out | right_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_32_read_out : '0;
  assign pe_32_left = (!(par_done_reg171_out | right_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg200_out | right_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg218_out | right_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg227_out | right_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_32_read_out : '0;
  assign pe_32_go = (!pe_32_done & (!(par_done_reg171_out | right_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg200_out | right_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg218_out | right_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg227_out | right_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_31_write_in = (pe_31_done & (!(par_done_reg133_out | right_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg170_out | right_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg199_out | right_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg217_out | right_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_31_right : '0;
  assign right_31_write_write_en = (pe_31_done & (!(par_done_reg133_out | right_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg170_out | right_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg199_out | right_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg217_out | right_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_31_read_in = (!(par_done_reg117_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg156_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg189_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg211_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_30_write_out : '0;
  assign left_31_read_write_en = (!(par_done_reg117_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg156_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg189_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg211_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_31_read_in = (!(par_done_reg105_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg144_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg179_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg205_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_21_write_out : '0;
  assign top_31_read_write_en = (!(par_done_reg105_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg144_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg179_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg205_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_31_top = (!(par_done_reg133_out | right_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg170_out | right_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg199_out | right_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg217_out | right_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_31_read_out : '0;
  assign pe_31_left = (!(par_done_reg133_out | right_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg170_out | right_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg199_out | right_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg217_out | right_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_31_read_out : '0;
  assign pe_31_go = (!pe_31_done & (!(par_done_reg133_out | right_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg170_out | right_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg199_out | right_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg217_out | right_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_30_write_in = (pe_30_done & (!(par_done_reg93_out | right_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | right_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg169_out | right_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg198_out | right_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_30_right : '0;
  assign right_30_write_write_en = (pe_30_done & (!(par_done_reg93_out | right_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | right_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg169_out | right_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg198_out | right_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_30_read_in = (!(par_done_reg77_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg155_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg188_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? l3_read_data : '0;
  assign left_30_read_write_en = (!(par_done_reg77_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg155_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg188_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_30_read_in = (!(par_done_reg67_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg104_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg143_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg178_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_20_write_out : '0;
  assign top_30_read_write_en = (!(par_done_reg67_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg104_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg143_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg178_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_30_top = (!(par_done_reg93_out | right_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | right_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg169_out | right_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg198_out | right_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_30_read_out : '0;
  assign pe_30_left = (!(par_done_reg93_out | right_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | right_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg169_out | right_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg198_out | right_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_30_read_out : '0;
  assign pe_30_go = (!pe_30_done & (!(par_done_reg93_out | right_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | right_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg169_out | right_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg198_out | right_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_23_write_in = (pe_23_done & (!(par_done_reg168_out | down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg197_out | down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg216_out | down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg226_out | down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_23_down : '0;
  assign down_23_write_write_en = (pe_23_done & (!(par_done_reg168_out | down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg197_out | down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg216_out | down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg226_out | down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_23_read_in = (!(par_done_reg154_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg187_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg210_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg223_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_22_write_out : '0;
  assign left_23_read_write_en = (!(par_done_reg154_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg187_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg210_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg223_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_23_read_in = (!(par_done_reg142_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg177_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg204_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg220_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_13_write_out : '0;
  assign top_23_read_write_en = (!(par_done_reg142_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg177_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg204_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg220_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_23_top = (!(par_done_reg168_out | down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg197_out | down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg216_out | down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg226_out | down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_23_read_out : '0;
  assign pe_23_left = (!(par_done_reg168_out | down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg197_out | down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg216_out | down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg226_out | down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_23_read_out : '0;
  assign pe_23_go = (!pe_23_done & (!(par_done_reg168_out | down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg197_out | down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg216_out | down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg226_out | down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_22_write_in = (pe_22_done & (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_22_down : '0;
  assign down_22_write_write_en = (pe_22_done & (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_22_write_in = (pe_22_done & (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_22_right : '0;
  assign right_22_write_write_en = (pe_22_done & (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_22_read_in = (!(par_done_reg115_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg153_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg186_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg209_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_21_write_out : '0;
  assign left_22_read_write_en = (!(par_done_reg115_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg153_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg186_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg209_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_22_read_in = (!(par_done_reg103_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg141_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg176_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg203_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_12_write_out : '0;
  assign top_22_read_write_en = (!(par_done_reg103_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg141_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg176_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg203_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_22_top = (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_22_read_out : '0;
  assign pe_22_left = (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_22_read_out : '0;
  assign pe_22_go = (!pe_22_done & (!(par_done_reg131_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg167_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg196_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg215_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_21_write_in = (pe_21_done & (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_21_down : '0;
  assign down_21_write_write_en = (pe_21_done & (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_21_write_in = (pe_21_done & (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_21_right : '0;
  assign right_21_write_write_en = (pe_21_done & (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_21_read_in = (!(par_done_reg76_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg114_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg152_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg185_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_20_write_out : '0;
  assign left_21_read_write_en = (!(par_done_reg76_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg114_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg152_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg185_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_21_read_in = (!(par_done_reg66_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg140_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg175_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_11_write_out : '0;
  assign top_21_read_write_en = (!(par_done_reg66_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg140_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg175_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_21_top = (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_21_read_out : '0;
  assign pe_21_left = (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_21_read_out : '0;
  assign pe_21_go = (!pe_21_done & (!(par_done_reg92_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg130_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg166_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg195_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_20_write_in = (pe_20_done & (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_20_down : '0;
  assign down_20_write_write_en = (pe_20_done & (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_20_write_in = (pe_20_done & (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_20_right : '0;
  assign right_20_write_write_en = (pe_20_done & (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_20_read_in = (!(par_done_reg43_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg75_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg113_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg151_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? l2_read_data : '0;
  assign left_20_read_write_en = (!(par_done_reg43_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg75_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg113_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg151_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_20_read_in = (!(par_done_reg37_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg65_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg101_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg139_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? down_10_write_out : '0;
  assign top_20_read_write_en = (!(par_done_reg37_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg65_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg101_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg139_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_20_top = (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_20_read_out : '0;
  assign pe_20_left = (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_20_read_out : '0;
  assign pe_20_go = (!pe_20_done & (!(par_done_reg57_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg91_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg129_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg165_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign down_13_write_in = (pe_13_done & (!(par_done_reg128_out | down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg164_out | down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg194_out | down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg214_out | down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_13_down : '0;
  assign down_13_write_write_en = (pe_13_done & (!(par_done_reg128_out | down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg164_out | down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg194_out | down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg214_out | down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_13_read_in = (!(par_done_reg112_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg150_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg184_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg208_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_12_write_out : '0;
  assign left_13_read_write_en = (!(par_done_reg112_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg150_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg184_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg208_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_13_read_in = (!(par_done_reg100_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg138_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg174_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg202_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_03_write_out : '0;
  assign top_13_read_write_en = (!(par_done_reg100_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg138_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg174_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg202_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_13_top = (!(par_done_reg128_out | down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg164_out | down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg194_out | down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg214_out | down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_13_read_out : '0;
  assign pe_13_left = (!(par_done_reg128_out | down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg164_out | down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg194_out | down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg214_out | down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_13_read_out : '0;
  assign pe_13_go = (!pe_13_done & (!(par_done_reg128_out | down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg164_out | down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg194_out | down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg214_out | down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_12_write_in = (pe_12_done & (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_12_down : '0;
  assign down_12_write_write_en = (pe_12_done & (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_12_write_in = (pe_12_done & (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_12_right : '0;
  assign right_12_write_write_en = (pe_12_done & (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_12_read_in = (!(par_done_reg74_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg111_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg149_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg183_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_11_write_out : '0;
  assign left_12_read_write_en = (!(par_done_reg74_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg111_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg149_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg183_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_12_read_in = (!(par_done_reg64_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg99_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg137_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg173_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_02_write_out : '0;
  assign top_12_read_write_en = (!(par_done_reg64_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg99_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg137_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg173_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_12_top = (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_12_read_out : '0;
  assign pe_12_left = (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_12_read_out : '0;
  assign pe_12_go = (!pe_12_done & (!(par_done_reg90_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg127_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg163_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg193_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_11_write_in = (pe_11_done & (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_11_down : '0;
  assign down_11_write_write_en = (pe_11_done & (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_11_write_in = (pe_11_done & (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_11_right : '0;
  assign right_11_write_write_en = (pe_11_done & (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_11_read_in = (!(par_done_reg42_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg73_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg110_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg148_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? right_10_write_out : '0;
  assign left_11_read_write_en = (!(par_done_reg42_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg73_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg110_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg148_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_11_read_in = (!(par_done_reg36_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg63_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg98_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg136_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? down_01_write_out : '0;
  assign top_11_read_write_en = (!(par_done_reg36_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg63_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg98_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg136_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_11_top = (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_11_read_out : '0;
  assign pe_11_left = (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_11_read_out : '0;
  assign pe_11_go = (!pe_11_done & (!(par_done_reg56_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg126_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg162_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign down_10_write_in = (pe_10_done & (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_10_down : '0;
  assign down_10_write_write_en = (pe_10_done & (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign right_10_write_in = (pe_10_done & (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_10_right : '0;
  assign right_10_write_write_en = (pe_10_done & (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign left_10_read_in = (!(par_done_reg22_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? l1_read_data : '0;
  assign left_10_read_write_en = (!(par_done_reg22_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign top_10_read_in = (!(par_done_reg19_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg35_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg97_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? down_00_write_out : '0;
  assign top_10_read_write_en = (!(par_done_reg19_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg35_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg97_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign pe_10_top = (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? top_10_read_out : '0;
  assign pe_10_left = (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? left_10_read_out : '0;
  assign pe_10_go = (!pe_10_done & (!(par_done_reg31_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg125_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign down_03_write_in = (pe_03_done & (!(par_done_reg87_out | down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg124_out | down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg161_out | down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg192_out | down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_03_down : '0;
  assign down_03_write_write_en = (pe_03_done & (!(par_done_reg87_out | down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg124_out | down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg161_out | down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg192_out | down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_03_read_in = (!(par_done_reg71_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg147_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg182_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_02_write_out : '0;
  assign left_03_read_write_en = (!(par_done_reg71_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg147_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg182_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_03_read_in = (!(par_done_reg61_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg96_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg135_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg172_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? t3_read_data : '0;
  assign top_03_read_write_en = (!(par_done_reg61_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg96_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg135_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg172_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_03_top = (!(par_done_reg87_out | down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg124_out | down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg161_out | down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg192_out | down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_03_read_out : '0;
  assign pe_03_left = (!(par_done_reg87_out | down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg124_out | down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg161_out | down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg192_out | down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_03_read_out : '0;
  assign pe_03_go = (!pe_03_done & (!(par_done_reg87_out | down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg124_out | down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg161_out | down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg192_out | down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_02_write_in = (pe_02_done & (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_02_down : '0;
  assign down_02_write_write_en = (pe_02_done & (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_02_write_in = (pe_02_done & (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_02_right : '0;
  assign right_02_write_write_en = (pe_02_done & (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_02_read_in = (!(par_done_reg40_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg146_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? right_01_write_out : '0;
  assign left_02_read_write_en = (!(par_done_reg40_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg146_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_02_read_in = (!(par_done_reg34_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg95_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg134_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? t2_read_data : '0;
  assign top_02_read_write_en = (!(par_done_reg34_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg95_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg134_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_02_top = (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_02_read_out : '0;
  assign pe_02_left = (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_02_read_out : '0;
  assign pe_02_go = (!pe_02_done & (!(par_done_reg54_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg123_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg160_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign down_01_write_in = (pe_01_done & (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_01_down : '0;
  assign down_01_write_write_en = (pe_01_done & (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign right_01_write_in = (pe_01_done & (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? pe_01_right : '0;
  assign right_01_write_write_en = (pe_01_done & (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign left_01_read_in = (!(par_done_reg21_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg69_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? right_00_write_out : '0;
  assign left_01_read_write_en = (!(par_done_reg21_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg69_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign top_01_read_in = (!(par_done_reg18_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg33_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg59_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg94_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? t1_read_data : '0;
  assign top_01_read_write_en = (!(par_done_reg18_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg33_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg59_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg94_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign pe_01_top = (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? top_01_read_out : '0;
  assign pe_01_left = (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? left_01_read_out : '0;
  assign pe_01_go = (!pe_01_done & (!(par_done_reg30_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg122_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go)) ? 1'd1 : '0;
  assign down_00_write_in = (pe_00_done & (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? pe_00_down : '0;
  assign down_00_write_write_en = (pe_00_done & (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign right_00_write_in = (pe_00_done & (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? pe_00_right : '0;
  assign right_00_write_write_en = (pe_00_done & (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign left_00_read_in = (!(par_done_reg11_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg20_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg38_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg68_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? l0_read_data : '0;
  assign left_00_read_write_en = (!(par_done_reg11_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg20_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg38_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg68_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign top_00_read_in = (!(par_done_reg10_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg17_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg32_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg58_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? t0_read_data : '0;
  assign top_00_read_write_en = (!(par_done_reg10_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg17_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg32_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg58_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign pe_00_top = (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? top_00_read_out : '0;
  assign pe_00_left = (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? left_00_read_out : '0;
  assign pe_00_go = (!pe_00_done & (!(par_done_reg16_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go)) ? 1'd1 : '0;
  assign l3_addr0 = (!(par_done_reg77_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg155_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg188_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? l3_idx_out : '0;
  assign l3_add_left = (!(par_done_reg51_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg121_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg159_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 3'd1 : '0;
  assign l3_add_right = (!(par_done_reg51_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg121_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg159_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? l3_idx_out : '0;
  assign l3_idx_in = (!(par_done_reg51_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg121_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg159_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? l3_add_out : (!(par_done_reg7_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l3_idx_write_en = (!(par_done_reg7_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg51_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg121_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg159_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign l2_addr0 = (!(par_done_reg43_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg75_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg113_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg151_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? l2_idx_out : '0;
  assign l2_add_left = (!(par_done_reg28_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg120_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 3'd1 : '0;
  assign l2_add_right = (!(par_done_reg28_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg120_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? l2_idx_out : '0;
  assign l2_idx_in = (!(par_done_reg28_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg120_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? l2_add_out : (!(par_done_reg6_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l2_idx_write_en = (!(par_done_reg6_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg28_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg120_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign l1_addr0 = (!(par_done_reg22_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? l1_idx_out : '0;
  assign l1_add_left = (!(par_done_reg15_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 3'd1 : '0;
  assign l1_add_right = (!(par_done_reg15_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? l1_idx_out : '0;
  assign l1_idx_in = (!(par_done_reg15_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? l1_add_out : (!(par_done_reg5_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l1_idx_write_en = (!(par_done_reg5_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg15_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg81_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign l0_addr0 = (!(par_done_reg11_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg20_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg38_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg68_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? l0_idx_out : '0;
  assign l0_add_left = (!(par_done_reg9_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg24_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 3'd1 : '0;
  assign l0_add_right = (!(par_done_reg9_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg24_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? l0_idx_out : '0;
  assign l0_idx_in = (!(par_done_reg9_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg24_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? l0_add_out : (!(par_done_reg4_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l0_idx_write_en = (!(par_done_reg4_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg9_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg24_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg45_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign t3_addr0 = (!(par_done_reg61_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg96_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg135_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg172_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? t3_idx_out : '0;
  assign t3_add_left = (!(par_done_reg48_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg119_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg158_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 3'd1 : '0;
  assign t3_add_right = (!(par_done_reg48_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg119_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg158_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? t3_idx_out : '0;
  assign t3_idx_in = (!(par_done_reg48_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg119_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg158_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? t3_add_out : (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t3_idx_write_en = (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg48_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg80_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg119_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg158_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign t2_addr0 = (!(par_done_reg34_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg60_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg95_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg134_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? t2_idx_out : '0;
  assign t2_add_left = (!(par_done_reg26_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg79_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg118_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 3'd1 : '0;
  assign t2_add_right = (!(par_done_reg26_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg79_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg118_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? t2_idx_out : '0;
  assign t2_idx_in = (!(par_done_reg26_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg79_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg118_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? t2_add_out : (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t2_idx_write_en = (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg26_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg47_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg79_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg118_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign t1_addr0 = (!(par_done_reg18_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg33_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg59_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg94_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go) ? t1_idx_out : '0;
  assign t1_add_left = (!(par_done_reg14_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg78_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 3'd1 : '0;
  assign t1_add_right = (!(par_done_reg14_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg78_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? t1_idx_out : '0;
  assign t1_idx_in = (!(par_done_reg14_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg78_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? t1_add_out : (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t1_idx_write_en = (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg14_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg25_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg46_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg78_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign t0_addr0 = (!(par_done_reg10_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg17_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg32_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg58_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go) ? t0_idx_out : '0;
  assign t0_add_left = (!(par_done_reg8_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 3'd1 : '0;
  assign t0_add_right = (!(par_done_reg8_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? t0_idx_out : '0;
  assign t0_idx_in = (!(par_done_reg8_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? t0_add_out : (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t0_idx_write_en = (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg8_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg23_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg44_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_reset0_in = par_reset0_out ? 1'd0 : (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_reset0_write_en = (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg0_in = par_reset0_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg0_write_en = (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg1_in = par_reset0_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg1_write_en = (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg2_in = par_reset0_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg2_write_en = (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg3_in = par_reset0_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg3_write_en = (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg4_in = par_reset0_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg4_write_en = (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg5_in = par_reset0_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg5_write_en = (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg6_in = par_reset0_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg6_write_en = (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg7_in = par_reset0_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg7_write_en = (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_reset1_in = par_reset1_out ? 1'd0 : (par_done_reg8_out & par_done_reg9_out & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_reset1_write_en = (par_done_reg8_out & par_done_reg9_out & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg8_in = par_reset1_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg8_write_en = (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg9_in = par_reset1_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg9_write_en = (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_reset2_in = par_reset2_out ? 1'd0 : (par_done_reg10_out & par_done_reg11_out & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_reset2_write_en = (par_done_reg10_out & par_done_reg11_out & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg10_in = par_reset2_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg10_write_en = (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg11_in = par_reset2_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg11_write_en = (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_reset3_in = par_reset3_out ? 1'd0 : (par_done_reg12_out & par_done_reg13_out & par_done_reg14_out & par_done_reg15_out & par_done_reg16_out & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_reset3_write_en = (par_done_reg12_out & par_done_reg13_out & par_done_reg14_out & par_done_reg15_out & par_done_reg16_out & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg12_in = par_reset3_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg12_write_en = (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg13_in = par_reset3_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg13_write_en = (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg14_in = par_reset3_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg14_write_en = (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg15_in = par_reset3_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg15_write_en = (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg16_in = par_reset3_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg16_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_reset4_in = par_reset4_out ? 1'd0 : (par_done_reg17_out & par_done_reg18_out & par_done_reg19_out & par_done_reg20_out & par_done_reg21_out & par_done_reg22_out & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_reset4_write_en = (par_done_reg17_out & par_done_reg18_out & par_done_reg19_out & par_done_reg20_out & par_done_reg21_out & par_done_reg22_out & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg17_in = par_reset4_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg17_write_en = (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg18_in = par_reset4_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg18_write_en = (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg19_in = par_reset4_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg19_write_en = (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg20_in = par_reset4_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg20_write_en = (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg21_in = par_reset4_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg21_write_en = (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg22_in = par_reset4_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg22_write_en = (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_reset5_in = par_reset5_out ? 1'd0 : (par_done_reg23_out & par_done_reg24_out & par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & par_done_reg31_out & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_reset5_write_en = (par_done_reg23_out & par_done_reg24_out & par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & par_done_reg31_out & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg23_in = par_reset5_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg23_write_en = (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg24_in = par_reset5_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg24_write_en = (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg25_in = par_reset5_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg25_write_en = (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg26_in = par_reset5_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg26_write_en = (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg27_in = par_reset5_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg27_write_en = (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg28_in = par_reset5_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg28_write_en = (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg29_in = par_reset5_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg29_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg30_in = par_reset5_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg30_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg31_in = par_reset5_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg31_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_reset6_in = par_reset6_out ? 1'd0 : (par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_reset6_write_en = (par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg32_in = par_reset6_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg32_write_en = (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg33_in = par_reset6_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg33_write_en = (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg34_in = par_reset6_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg34_write_en = (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg35_in = par_reset6_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg35_write_en = (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg36_in = par_reset6_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg36_write_en = (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg37_in = par_reset6_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg37_write_en = (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg38_in = par_reset6_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg38_write_en = (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg39_in = par_reset6_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg39_write_en = (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg40_in = par_reset6_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg40_write_en = (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg41_in = par_reset6_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg41_write_en = (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg42_in = par_reset6_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg42_write_en = (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg43_in = par_reset6_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg43_write_en = (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_reset7_in = par_reset7_out ? 1'd0 : (par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_reset7_write_en = (par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg44_in = par_reset7_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg44_write_en = (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg45_in = par_reset7_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg45_write_en = (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg46_in = par_reset7_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg46_write_en = (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg47_in = par_reset7_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg47_write_en = (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg48_in = par_reset7_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg48_write_en = (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg49_in = par_reset7_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg49_write_en = (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg50_in = par_reset7_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg50_write_en = (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg51_in = par_reset7_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg51_write_en = (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg52_in = par_reset7_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg52_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg53_in = par_reset7_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg53_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg54_in = par_reset7_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg54_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg55_in = par_reset7_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg55_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg56_in = par_reset7_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg56_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg57_in = par_reset7_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg57_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_reset8_in = par_reset8_out ? 1'd0 : (par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_reset8_write_en = (par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg58_in = par_reset8_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg58_write_en = (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg59_in = par_reset8_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg59_write_en = (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg60_in = par_reset8_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg60_write_en = (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg61_in = par_reset8_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg61_write_en = (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg62_in = par_reset8_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg62_write_en = (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg63_in = par_reset8_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg63_write_en = (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg64_in = par_reset8_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg64_write_en = (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg65_in = par_reset8_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg65_write_en = (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg66_in = par_reset8_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg66_write_en = (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg67_in = par_reset8_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg67_write_en = (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg68_in = par_reset8_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg68_write_en = (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg69_in = par_reset8_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg69_write_en = (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg70_in = par_reset8_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg70_write_en = (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg71_in = par_reset8_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg71_write_en = (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg72_in = par_reset8_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg72_write_en = (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg73_in = par_reset8_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg73_write_en = (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg74_in = par_reset8_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg74_write_en = (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg75_in = par_reset8_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg75_write_en = (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg76_in = par_reset8_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg76_write_en = (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg77_in = par_reset8_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg77_write_en = (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_reset9_in = par_reset9_out ? 1'd0 : (par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_reset9_write_en = (par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg78_in = par_reset9_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg78_write_en = (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg79_in = par_reset9_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg79_write_en = (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg80_in = par_reset9_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg80_write_en = (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg81_in = par_reset9_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg81_write_en = (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg82_in = par_reset9_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg82_write_en = (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg83_in = par_reset9_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg83_write_en = (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg84_in = par_reset9_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg84_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg85_in = par_reset9_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg85_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg86_in = par_reset9_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg86_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg87_in = par_reset9_out ? 1'd0 : (down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg87_write_en = (down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg88_in = par_reset9_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg88_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg89_in = par_reset9_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg89_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg90_in = par_reset9_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg90_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg91_in = par_reset9_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg91_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg92_in = par_reset9_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg92_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg93_in = par_reset9_out ? 1'd0 : (right_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg93_write_en = (right_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_reset10_in = par_reset10_out ? 1'd0 : (par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_reset10_write_en = (par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg94_in = par_reset10_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg94_write_en = (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg95_in = par_reset10_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg95_write_en = (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg96_in = par_reset10_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg96_write_en = (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg97_in = par_reset10_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg97_write_en = (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg98_in = par_reset10_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg98_write_en = (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg99_in = par_reset10_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg99_write_en = (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg100_in = par_reset10_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg100_write_en = (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg101_in = par_reset10_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg101_write_en = (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg102_in = par_reset10_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg102_write_en = (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg103_in = par_reset10_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg103_write_en = (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg104_in = par_reset10_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg104_write_en = (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg105_in = par_reset10_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg105_write_en = (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg106_in = par_reset10_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg106_write_en = (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg107_in = par_reset10_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg107_write_en = (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg108_in = par_reset10_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg108_write_en = (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg109_in = par_reset10_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg109_write_en = (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg110_in = par_reset10_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg110_write_en = (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg111_in = par_reset10_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg111_write_en = (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg112_in = par_reset10_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg112_write_en = (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg113_in = par_reset10_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg113_write_en = (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg114_in = par_reset10_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg114_write_en = (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg115_in = par_reset10_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg115_write_en = (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg116_in = par_reset10_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg116_write_en = (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg117_in = par_reset10_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg117_write_en = (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_reset11_in = par_reset11_out ? 1'd0 : (par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & par_done_reg130_out & par_done_reg131_out & par_done_reg132_out & par_done_reg133_out & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_reset11_write_en = (par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & par_done_reg130_out & par_done_reg131_out & par_done_reg132_out & par_done_reg133_out & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg118_in = par_reset11_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg118_write_en = (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg119_in = par_reset11_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg119_write_en = (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg120_in = par_reset11_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg120_write_en = (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg121_in = par_reset11_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg121_write_en = (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg122_in = par_reset11_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg122_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg123_in = par_reset11_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg123_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg124_in = par_reset11_out ? 1'd0 : (down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg124_write_en = (down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg125_in = par_reset11_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg125_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg126_in = par_reset11_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg126_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg127_in = par_reset11_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg127_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg128_in = par_reset11_out ? 1'd0 : (down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg128_write_en = (down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg129_in = par_reset11_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg129_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg130_in = par_reset11_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg130_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg131_in = par_reset11_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg131_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg132_in = par_reset11_out ? 1'd0 : (right_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg132_write_en = (right_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg133_in = par_reset11_out ? 1'd0 : (right_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg133_write_en = (right_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_reset12_in = par_reset12_out ? 1'd0 : (par_done_reg134_out & par_done_reg135_out & par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_reset12_write_en = (par_done_reg134_out & par_done_reg135_out & par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg134_in = par_reset12_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg134_write_en = (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg135_in = par_reset12_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg135_write_en = (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg136_in = par_reset12_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg136_write_en = (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg137_in = par_reset12_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg137_write_en = (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg138_in = par_reset12_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg138_write_en = (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg139_in = par_reset12_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg139_write_en = (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg140_in = par_reset12_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg140_write_en = (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg141_in = par_reset12_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg141_write_en = (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg142_in = par_reset12_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg142_write_en = (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg143_in = par_reset12_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg143_write_en = (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg144_in = par_reset12_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg144_write_en = (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg145_in = par_reset12_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg145_write_en = (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg146_in = par_reset12_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg146_write_en = (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg147_in = par_reset12_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg147_write_en = (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg148_in = par_reset12_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg148_write_en = (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg149_in = par_reset12_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg149_write_en = (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg150_in = par_reset12_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg150_write_en = (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg151_in = par_reset12_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg151_write_en = (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg152_in = par_reset12_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg152_write_en = (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg153_in = par_reset12_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg153_write_en = (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg154_in = par_reset12_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg154_write_en = (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg155_in = par_reset12_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg155_write_en = (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg156_in = par_reset12_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg156_write_en = (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg157_in = par_reset12_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg157_write_en = (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_reset13_in = par_reset13_out ? 1'd0 : (par_done_reg158_out & par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_reset13_write_en = (par_done_reg158_out & par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg158_in = par_reset13_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg158_write_en = (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg159_in = par_reset13_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg159_write_en = (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg160_in = par_reset13_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg160_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg161_in = par_reset13_out ? 1'd0 : (down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg161_write_en = (down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg162_in = par_reset13_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg162_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg163_in = par_reset13_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg163_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg164_in = par_reset13_out ? 1'd0 : (down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg164_write_en = (down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg165_in = par_reset13_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg165_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg166_in = par_reset13_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg166_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg167_in = par_reset13_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg167_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg168_in = par_reset13_out ? 1'd0 : (down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg168_write_en = (down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg169_in = par_reset13_out ? 1'd0 : (right_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg169_write_en = (right_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg170_in = par_reset13_out ? 1'd0 : (right_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg170_write_en = (right_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg171_in = par_reset13_out ? 1'd0 : (right_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg171_write_en = (right_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_reset14_in = par_reset14_out ? 1'd0 : (par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_reset14_write_en = (par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg172_in = par_reset14_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg172_write_en = (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg173_in = par_reset14_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg173_write_en = (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg174_in = par_reset14_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg174_write_en = (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg175_in = par_reset14_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg175_write_en = (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg176_in = par_reset14_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg176_write_en = (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg177_in = par_reset14_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg177_write_en = (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg178_in = par_reset14_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg178_write_en = (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg179_in = par_reset14_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg179_write_en = (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg180_in = par_reset14_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg180_write_en = (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg181_in = par_reset14_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg181_write_en = (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg182_in = par_reset14_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg182_write_en = (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg183_in = par_reset14_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg183_write_en = (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg184_in = par_reset14_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg184_write_en = (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg185_in = par_reset14_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg185_write_en = (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg186_in = par_reset14_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg186_write_en = (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg187_in = par_reset14_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg187_write_en = (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg188_in = par_reset14_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg188_write_en = (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg189_in = par_reset14_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg189_write_en = (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg190_in = par_reset14_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg190_write_en = (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg191_in = par_reset14_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg191_write_en = (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_reset15_in = par_reset15_out ? 1'd0 : (par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & par_done_reg201_out & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_reset15_write_en = (par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & par_done_reg201_out & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg192_in = par_reset15_out ? 1'd0 : (down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg192_write_en = (down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg193_in = par_reset15_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg193_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg194_in = par_reset15_out ? 1'd0 : (down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg194_write_en = (down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg195_in = par_reset15_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg195_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg196_in = par_reset15_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg196_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg197_in = par_reset15_out ? 1'd0 : (down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg197_write_en = (down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg198_in = par_reset15_out ? 1'd0 : (right_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg198_write_en = (right_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg199_in = par_reset15_out ? 1'd0 : (right_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg199_write_en = (right_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg200_in = par_reset15_out ? 1'd0 : (right_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg200_write_en = (right_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg201_in = par_reset15_out ? 1'd0 : (pe_33_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg201_write_en = (pe_33_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_reset16_in = par_reset16_out ? 1'd0 : (par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & par_done_reg213_out & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_reset16_write_en = (par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & par_done_reg213_out & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg202_in = par_reset16_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg202_write_en = (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg203_in = par_reset16_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg203_write_en = (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg204_in = par_reset16_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg204_write_en = (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg205_in = par_reset16_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg205_write_en = (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg206_in = par_reset16_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg206_write_en = (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg207_in = par_reset16_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg207_write_en = (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg208_in = par_reset16_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg208_write_en = (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg209_in = par_reset16_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg209_write_en = (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg210_in = par_reset16_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg210_write_en = (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg211_in = par_reset16_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg211_write_en = (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg212_in = par_reset16_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg212_write_en = (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg213_in = par_reset16_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg213_write_en = (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_reset17_in = par_reset17_out ? 1'd0 : (par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_reset17_write_en = (par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg214_in = par_reset17_out ? 1'd0 : (down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg214_write_en = (down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg215_in = par_reset17_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg215_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg216_in = par_reset17_out ? 1'd0 : (down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg216_write_en = (down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg217_in = par_reset17_out ? 1'd0 : (right_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg217_write_en = (right_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg218_in = par_reset17_out ? 1'd0 : (right_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg218_write_en = (right_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg219_in = par_reset17_out ? 1'd0 : (pe_33_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg219_write_en = (pe_33_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_reset18_in = par_reset18_out ? 1'd0 : (par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_reset18_write_en = (par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg220_in = par_reset18_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg220_write_en = (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg221_in = par_reset18_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg221_write_en = (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg222_in = par_reset18_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg222_write_en = (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg223_in = par_reset18_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg223_write_en = (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg224_in = par_reset18_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg224_write_en = (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg225_in = par_reset18_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg225_write_en = (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_reset19_in = par_reset19_out ? 1'd0 : (par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_reset19_write_en = (par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg226_in = par_reset19_out ? 1'd0 : (down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg226_write_en = (down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg227_in = par_reset19_out ? 1'd0 : (right_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg227_write_en = (right_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg228_in = par_reset19_out ? 1'd0 : (pe_33_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg228_write_en = (pe_33_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_reset20_in = par_reset20_out ? 1'd0 : (par_done_reg229_out & par_done_reg230_out & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_reset20_write_en = (par_done_reg229_out & par_done_reg230_out & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg229_in = par_reset20_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg229_write_en = (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg230_in = par_reset20_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg230_write_en = (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_reset21_in = par_reset21_out ? 1'd0 : (par_done_reg231_out & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_reset21_write_en = (par_done_reg231_out & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg231_in = par_reset21_out ? 1'd0 : (pe_33_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg231_write_en = (pe_33_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd1 & par_reset1_out & go) ? 32'd2 : (fsm0_out == 32'd0 & par_reset0_out & go) ? 32'd1 : (fsm0_out == 32'd38) ? 32'd0 : (fsm0_out == 32'd37 & out_mem_done & go) ? 32'd38 : (fsm0_out == 32'd36 & out_mem_done & go) ? 32'd37 : (fsm0_out == 32'd35 & out_mem_done & go) ? 32'd36 : (fsm0_out == 32'd34 & out_mem_done & go) ? 32'd35 : (fsm0_out == 32'd33 & out_mem_done & go) ? 32'd34 : (fsm0_out == 32'd32 & out_mem_done & go) ? 32'd33 : (fsm0_out == 32'd31 & out_mem_done & go) ? 32'd32 : (fsm0_out == 32'd30 & out_mem_done & go) ? 32'd31 : (fsm0_out == 32'd29 & out_mem_done & go) ? 32'd30 : (fsm0_out == 32'd28 & out_mem_done & go) ? 32'd29 : (fsm0_out == 32'd27 & out_mem_done & go) ? 32'd28 : (fsm0_out == 32'd26 & out_mem_done & go) ? 32'd27 : (fsm0_out == 32'd25 & out_mem_done & go) ? 32'd26 : (fsm0_out == 32'd24 & out_mem_done & go) ? 32'd25 : (fsm0_out == 32'd23 & out_mem_done & go) ? 32'd24 : (fsm0_out == 32'd22 & out_mem_done & go) ? 32'd23 : (fsm0_out == 32'd21 & par_reset21_out & go) ? 32'd22 : (fsm0_out == 32'd20 & par_reset20_out & go) ? 32'd21 : (fsm0_out == 32'd19 & par_reset19_out & go) ? 32'd20 : (fsm0_out == 32'd18 & par_reset18_out & go) ? 32'd19 : (fsm0_out == 32'd17 & par_reset17_out & go) ? 32'd18 : (fsm0_out == 32'd16 & par_reset16_out & go) ? 32'd17 : (fsm0_out == 32'd15 & par_reset15_out & go) ? 32'd16 : (fsm0_out == 32'd14 & par_reset14_out & go) ? 32'd15 : (fsm0_out == 32'd13 & par_reset13_out & go) ? 32'd14 : (fsm0_out == 32'd12 & par_reset12_out & go) ? 32'd13 : (fsm0_out == 32'd11 & par_reset11_out & go) ? 32'd12 : (fsm0_out == 32'd10 & par_reset10_out & go) ? 32'd11 : (fsm0_out == 32'd9 & par_reset9_out & go) ? 32'd10 : (fsm0_out == 32'd8 & par_reset8_out & go) ? 32'd9 : (fsm0_out == 32'd7 & par_reset7_out & go) ? 32'd8 : (fsm0_out == 32'd6 & par_reset6_out & go) ? 32'd7 : (fsm0_out == 32'd5 & par_reset5_out & go) ? 32'd6 : (fsm0_out == 32'd4 & par_reset4_out & go) ? 32'd5 : (fsm0_out == 32'd3 & par_reset3_out & go) ? 32'd4 : (fsm0_out == 32'd2 & par_reset2_out & go) ? 32'd3 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & par_reset0_out & go | fsm0_out == 32'd1 & par_reset1_out & go | fsm0_out == 32'd2 & par_reset2_out & go | fsm0_out == 32'd3 & par_reset3_out & go | fsm0_out == 32'd4 & par_reset4_out & go | fsm0_out == 32'd5 & par_reset5_out & go | fsm0_out == 32'd6 & par_reset6_out & go | fsm0_out == 32'd7 & par_reset7_out & go | fsm0_out == 32'd8 & par_reset8_out & go | fsm0_out == 32'd9 & par_reset9_out & go | fsm0_out == 32'd10 & par_reset10_out & go | fsm0_out == 32'd11 & par_reset11_out & go | fsm0_out == 32'd12 & par_reset12_out & go | fsm0_out == 32'd13 & par_reset13_out & go | fsm0_out == 32'd14 & par_reset14_out & go | fsm0_out == 32'd15 & par_reset15_out & go | fsm0_out == 32'd16 & par_reset16_out & go | fsm0_out == 32'd17 & par_reset17_out & go | fsm0_out == 32'd18 & par_reset18_out & go | fsm0_out == 32'd19 & par_reset19_out & go | fsm0_out == 32'd20 & par_reset20_out & go | fsm0_out == 32'd21 & par_reset21_out & go | fsm0_out == 32'd22 & out_mem_done & go | fsm0_out == 32'd23 & out_mem_done & go | fsm0_out == 32'd24 & out_mem_done & go | fsm0_out == 32'd25 & out_mem_done & go | fsm0_out == 32'd26 & out_mem_done & go | fsm0_out == 32'd27 & out_mem_done & go | fsm0_out == 32'd28 & out_mem_done & go | fsm0_out == 32'd29 & out_mem_done & go | fsm0_out == 32'd30 & out_mem_done & go | fsm0_out == 32'd31 & out_mem_done & go | fsm0_out == 32'd32 & out_mem_done & go | fsm0_out == 32'd33 & out_mem_done & go | fsm0_out == 32'd34 & out_mem_done & go | fsm0_out == 32'd35 & out_mem_done & go | fsm0_out == 32'd36 & out_mem_done & go | fsm0_out == 32'd37 & out_mem_done & go | fsm0_out == 32'd38) ? 1'd1 : '0;
endmodule // end main