/* verilator lint_off WIDTH */
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule

module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule

module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

// Component Signature
module mac_pe (
      input wire [31:0] top,
      input wire [31:0] left,
      input wire go,
      input wire clk,
      output wire [31:0] down,
      output wire [31:0] right,
      output wire [31:0] out,
      output wire done
  );
  
  // Structure wire declarations
  wire [31:0] mul_left;
  wire [31:0] mul_right;
  wire mul_go;
  wire mul_clk;
  wire [31:0] mul_out;
  wire mul_done;
  wire [31:0] add_left;
  wire [31:0] add_right;
  wire [31:0] add_out;
  wire [31:0] mul_reg_in;
  wire mul_reg_write_en;
  wire mul_reg_clk;
  wire [31:0] mul_reg_out;
  wire mul_reg_done;
  wire [31:0] acc_in;
  wire acc_write_en;
  wire acc_clk;
  wire [31:0] acc_out;
  wire acc_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_mult_pipe #(32) mul (
      .left(mul_left),
      .right(mul_right),
      .go(mul_go),
      .clk(clk),
      .out(mul_out),
      .done(mul_done)
  );
  
  std_add #(32) add (
      .left(add_left),
      .right(add_right),
      .out(add_out)
  );
  
  std_reg #(32) mul_reg (
      .in(mul_reg_in),
      .write_en(mul_reg_write_en),
      .clk(clk),
      .out(mul_reg_out),
      .done(mul_reg_done)
  );
  
  std_reg #(32) acc (
      .in(acc_in),
      .write_en(acc_write_en),
      .clk(clk),
      .out(acc_out),
      .done(acc_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign down = top;
  assign right = left;
  assign out = acc_out;
  assign done = (fsm0_out == 32'd2) ? 1'd1 : '0;
  assign mul_left = (fsm0_out == 32'd0 & !mul_reg_done & go) ? top : '0;
  assign mul_right = (fsm0_out == 32'd0 & !mul_reg_done & go) ? left : '0;
  assign mul_go = (!mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign add_left = (fsm0_out == 32'd1 & !acc_done & go) ? acc_out : '0;
  assign add_right = (fsm0_out == 32'd1 & !acc_done & go) ? mul_reg_out : '0;
  assign mul_reg_in = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? mul_out : '0;
  assign mul_reg_write_en = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign acc_in = (fsm0_out == 32'd1 & !acc_done & go) ? add_out : '0;
  assign acc_write_en = (fsm0_out == 32'd1 & !acc_done & go) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd1 & acc_done & go) ? 32'd2 : (fsm0_out == 32'd0 & mul_reg_done & go) ? 32'd1 : (fsm0_out == 32'd2) ? 32'd0 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & mul_reg_done & go | fsm0_out == 32'd1 & acc_done & go | fsm0_out == 32'd2) ? 1'd1 : '0;
endmodule // end mac_pe
// Component Signature
module main (
      input wire go,
      input wire clk,
      input wire [31:0] out_mem_read_data,
      input wire out_mem_done,
      output wire done,
      output wire [2:0] out_mem_addr0,
      output wire [2:0] out_mem_addr1,
      output wire [31:0] out_mem_write_data,
      output wire out_mem_write_en
  );
  
  // Structure wire declarations
  wire [31:0] left_55_read_in;
  wire left_55_read_write_en;
  wire left_55_read_clk;
  wire [31:0] left_55_read_out;
  wire left_55_read_done;
  wire [31:0] top_55_read_in;
  wire top_55_read_write_en;
  wire top_55_read_clk;
  wire [31:0] top_55_read_out;
  wire top_55_read_done;
  wire [31:0] pe_55_top;
  wire [31:0] pe_55_left;
  wire pe_55_go;
  wire pe_55_clk;
  wire [31:0] pe_55_down;
  wire [31:0] pe_55_right;
  wire [31:0] pe_55_out;
  wire pe_55_done;
  wire [31:0] right_54_write_in;
  wire right_54_write_write_en;
  wire right_54_write_clk;
  wire [31:0] right_54_write_out;
  wire right_54_write_done;
  wire [31:0] left_54_read_in;
  wire left_54_read_write_en;
  wire left_54_read_clk;
  wire [31:0] left_54_read_out;
  wire left_54_read_done;
  wire [31:0] top_54_read_in;
  wire top_54_read_write_en;
  wire top_54_read_clk;
  wire [31:0] top_54_read_out;
  wire top_54_read_done;
  wire [31:0] pe_54_top;
  wire [31:0] pe_54_left;
  wire pe_54_go;
  wire pe_54_clk;
  wire [31:0] pe_54_down;
  wire [31:0] pe_54_right;
  wire [31:0] pe_54_out;
  wire pe_54_done;
  wire [31:0] right_53_write_in;
  wire right_53_write_write_en;
  wire right_53_write_clk;
  wire [31:0] right_53_write_out;
  wire right_53_write_done;
  wire [31:0] left_53_read_in;
  wire left_53_read_write_en;
  wire left_53_read_clk;
  wire [31:0] left_53_read_out;
  wire left_53_read_done;
  wire [31:0] top_53_read_in;
  wire top_53_read_write_en;
  wire top_53_read_clk;
  wire [31:0] top_53_read_out;
  wire top_53_read_done;
  wire [31:0] pe_53_top;
  wire [31:0] pe_53_left;
  wire pe_53_go;
  wire pe_53_clk;
  wire [31:0] pe_53_down;
  wire [31:0] pe_53_right;
  wire [31:0] pe_53_out;
  wire pe_53_done;
  wire [31:0] right_52_write_in;
  wire right_52_write_write_en;
  wire right_52_write_clk;
  wire [31:0] right_52_write_out;
  wire right_52_write_done;
  wire [31:0] left_52_read_in;
  wire left_52_read_write_en;
  wire left_52_read_clk;
  wire [31:0] left_52_read_out;
  wire left_52_read_done;
  wire [31:0] top_52_read_in;
  wire top_52_read_write_en;
  wire top_52_read_clk;
  wire [31:0] top_52_read_out;
  wire top_52_read_done;
  wire [31:0] pe_52_top;
  wire [31:0] pe_52_left;
  wire pe_52_go;
  wire pe_52_clk;
  wire [31:0] pe_52_down;
  wire [31:0] pe_52_right;
  wire [31:0] pe_52_out;
  wire pe_52_done;
  wire [31:0] right_51_write_in;
  wire right_51_write_write_en;
  wire right_51_write_clk;
  wire [31:0] right_51_write_out;
  wire right_51_write_done;
  wire [31:0] left_51_read_in;
  wire left_51_read_write_en;
  wire left_51_read_clk;
  wire [31:0] left_51_read_out;
  wire left_51_read_done;
  wire [31:0] top_51_read_in;
  wire top_51_read_write_en;
  wire top_51_read_clk;
  wire [31:0] top_51_read_out;
  wire top_51_read_done;
  wire [31:0] pe_51_top;
  wire [31:0] pe_51_left;
  wire pe_51_go;
  wire pe_51_clk;
  wire [31:0] pe_51_down;
  wire [31:0] pe_51_right;
  wire [31:0] pe_51_out;
  wire pe_51_done;
  wire [31:0] right_50_write_in;
  wire right_50_write_write_en;
  wire right_50_write_clk;
  wire [31:0] right_50_write_out;
  wire right_50_write_done;
  wire [31:0] left_50_read_in;
  wire left_50_read_write_en;
  wire left_50_read_clk;
  wire [31:0] left_50_read_out;
  wire left_50_read_done;
  wire [31:0] top_50_read_in;
  wire top_50_read_write_en;
  wire top_50_read_clk;
  wire [31:0] top_50_read_out;
  wire top_50_read_done;
  wire [31:0] pe_50_top;
  wire [31:0] pe_50_left;
  wire pe_50_go;
  wire pe_50_clk;
  wire [31:0] pe_50_down;
  wire [31:0] pe_50_right;
  wire [31:0] pe_50_out;
  wire pe_50_done;
  wire [31:0] down_45_write_in;
  wire down_45_write_write_en;
  wire down_45_write_clk;
  wire [31:0] down_45_write_out;
  wire down_45_write_done;
  wire [31:0] left_45_read_in;
  wire left_45_read_write_en;
  wire left_45_read_clk;
  wire [31:0] left_45_read_out;
  wire left_45_read_done;
  wire [31:0] top_45_read_in;
  wire top_45_read_write_en;
  wire top_45_read_clk;
  wire [31:0] top_45_read_out;
  wire top_45_read_done;
  wire [31:0] pe_45_top;
  wire [31:0] pe_45_left;
  wire pe_45_go;
  wire pe_45_clk;
  wire [31:0] pe_45_down;
  wire [31:0] pe_45_right;
  wire [31:0] pe_45_out;
  wire pe_45_done;
  wire [31:0] down_44_write_in;
  wire down_44_write_write_en;
  wire down_44_write_clk;
  wire [31:0] down_44_write_out;
  wire down_44_write_done;
  wire [31:0] right_44_write_in;
  wire right_44_write_write_en;
  wire right_44_write_clk;
  wire [31:0] right_44_write_out;
  wire right_44_write_done;
  wire [31:0] left_44_read_in;
  wire left_44_read_write_en;
  wire left_44_read_clk;
  wire [31:0] left_44_read_out;
  wire left_44_read_done;
  wire [31:0] top_44_read_in;
  wire top_44_read_write_en;
  wire top_44_read_clk;
  wire [31:0] top_44_read_out;
  wire top_44_read_done;
  wire [31:0] pe_44_top;
  wire [31:0] pe_44_left;
  wire pe_44_go;
  wire pe_44_clk;
  wire [31:0] pe_44_down;
  wire [31:0] pe_44_right;
  wire [31:0] pe_44_out;
  wire pe_44_done;
  wire [31:0] down_43_write_in;
  wire down_43_write_write_en;
  wire down_43_write_clk;
  wire [31:0] down_43_write_out;
  wire down_43_write_done;
  wire [31:0] right_43_write_in;
  wire right_43_write_write_en;
  wire right_43_write_clk;
  wire [31:0] right_43_write_out;
  wire right_43_write_done;
  wire [31:0] left_43_read_in;
  wire left_43_read_write_en;
  wire left_43_read_clk;
  wire [31:0] left_43_read_out;
  wire left_43_read_done;
  wire [31:0] top_43_read_in;
  wire top_43_read_write_en;
  wire top_43_read_clk;
  wire [31:0] top_43_read_out;
  wire top_43_read_done;
  wire [31:0] pe_43_top;
  wire [31:0] pe_43_left;
  wire pe_43_go;
  wire pe_43_clk;
  wire [31:0] pe_43_down;
  wire [31:0] pe_43_right;
  wire [31:0] pe_43_out;
  wire pe_43_done;
  wire [31:0] down_42_write_in;
  wire down_42_write_write_en;
  wire down_42_write_clk;
  wire [31:0] down_42_write_out;
  wire down_42_write_done;
  wire [31:0] right_42_write_in;
  wire right_42_write_write_en;
  wire right_42_write_clk;
  wire [31:0] right_42_write_out;
  wire right_42_write_done;
  wire [31:0] left_42_read_in;
  wire left_42_read_write_en;
  wire left_42_read_clk;
  wire [31:0] left_42_read_out;
  wire left_42_read_done;
  wire [31:0] top_42_read_in;
  wire top_42_read_write_en;
  wire top_42_read_clk;
  wire [31:0] top_42_read_out;
  wire top_42_read_done;
  wire [31:0] pe_42_top;
  wire [31:0] pe_42_left;
  wire pe_42_go;
  wire pe_42_clk;
  wire [31:0] pe_42_down;
  wire [31:0] pe_42_right;
  wire [31:0] pe_42_out;
  wire pe_42_done;
  wire [31:0] down_41_write_in;
  wire down_41_write_write_en;
  wire down_41_write_clk;
  wire [31:0] down_41_write_out;
  wire down_41_write_done;
  wire [31:0] right_41_write_in;
  wire right_41_write_write_en;
  wire right_41_write_clk;
  wire [31:0] right_41_write_out;
  wire right_41_write_done;
  wire [31:0] left_41_read_in;
  wire left_41_read_write_en;
  wire left_41_read_clk;
  wire [31:0] left_41_read_out;
  wire left_41_read_done;
  wire [31:0] top_41_read_in;
  wire top_41_read_write_en;
  wire top_41_read_clk;
  wire [31:0] top_41_read_out;
  wire top_41_read_done;
  wire [31:0] pe_41_top;
  wire [31:0] pe_41_left;
  wire pe_41_go;
  wire pe_41_clk;
  wire [31:0] pe_41_down;
  wire [31:0] pe_41_right;
  wire [31:0] pe_41_out;
  wire pe_41_done;
  wire [31:0] down_40_write_in;
  wire down_40_write_write_en;
  wire down_40_write_clk;
  wire [31:0] down_40_write_out;
  wire down_40_write_done;
  wire [31:0] right_40_write_in;
  wire right_40_write_write_en;
  wire right_40_write_clk;
  wire [31:0] right_40_write_out;
  wire right_40_write_done;
  wire [31:0] left_40_read_in;
  wire left_40_read_write_en;
  wire left_40_read_clk;
  wire [31:0] left_40_read_out;
  wire left_40_read_done;
  wire [31:0] top_40_read_in;
  wire top_40_read_write_en;
  wire top_40_read_clk;
  wire [31:0] top_40_read_out;
  wire top_40_read_done;
  wire [31:0] pe_40_top;
  wire [31:0] pe_40_left;
  wire pe_40_go;
  wire pe_40_clk;
  wire [31:0] pe_40_down;
  wire [31:0] pe_40_right;
  wire [31:0] pe_40_out;
  wire pe_40_done;
  wire [31:0] down_35_write_in;
  wire down_35_write_write_en;
  wire down_35_write_clk;
  wire [31:0] down_35_write_out;
  wire down_35_write_done;
  wire [31:0] left_35_read_in;
  wire left_35_read_write_en;
  wire left_35_read_clk;
  wire [31:0] left_35_read_out;
  wire left_35_read_done;
  wire [31:0] top_35_read_in;
  wire top_35_read_write_en;
  wire top_35_read_clk;
  wire [31:0] top_35_read_out;
  wire top_35_read_done;
  wire [31:0] pe_35_top;
  wire [31:0] pe_35_left;
  wire pe_35_go;
  wire pe_35_clk;
  wire [31:0] pe_35_down;
  wire [31:0] pe_35_right;
  wire [31:0] pe_35_out;
  wire pe_35_done;
  wire [31:0] down_34_write_in;
  wire down_34_write_write_en;
  wire down_34_write_clk;
  wire [31:0] down_34_write_out;
  wire down_34_write_done;
  wire [31:0] right_34_write_in;
  wire right_34_write_write_en;
  wire right_34_write_clk;
  wire [31:0] right_34_write_out;
  wire right_34_write_done;
  wire [31:0] left_34_read_in;
  wire left_34_read_write_en;
  wire left_34_read_clk;
  wire [31:0] left_34_read_out;
  wire left_34_read_done;
  wire [31:0] top_34_read_in;
  wire top_34_read_write_en;
  wire top_34_read_clk;
  wire [31:0] top_34_read_out;
  wire top_34_read_done;
  wire [31:0] pe_34_top;
  wire [31:0] pe_34_left;
  wire pe_34_go;
  wire pe_34_clk;
  wire [31:0] pe_34_down;
  wire [31:0] pe_34_right;
  wire [31:0] pe_34_out;
  wire pe_34_done;
  wire [31:0] down_33_write_in;
  wire down_33_write_write_en;
  wire down_33_write_clk;
  wire [31:0] down_33_write_out;
  wire down_33_write_done;
  wire [31:0] right_33_write_in;
  wire right_33_write_write_en;
  wire right_33_write_clk;
  wire [31:0] right_33_write_out;
  wire right_33_write_done;
  wire [31:0] left_33_read_in;
  wire left_33_read_write_en;
  wire left_33_read_clk;
  wire [31:0] left_33_read_out;
  wire left_33_read_done;
  wire [31:0] top_33_read_in;
  wire top_33_read_write_en;
  wire top_33_read_clk;
  wire [31:0] top_33_read_out;
  wire top_33_read_done;
  wire [31:0] pe_33_top;
  wire [31:0] pe_33_left;
  wire pe_33_go;
  wire pe_33_clk;
  wire [31:0] pe_33_down;
  wire [31:0] pe_33_right;
  wire [31:0] pe_33_out;
  wire pe_33_done;
  wire [31:0] down_32_write_in;
  wire down_32_write_write_en;
  wire down_32_write_clk;
  wire [31:0] down_32_write_out;
  wire down_32_write_done;
  wire [31:0] right_32_write_in;
  wire right_32_write_write_en;
  wire right_32_write_clk;
  wire [31:0] right_32_write_out;
  wire right_32_write_done;
  wire [31:0] left_32_read_in;
  wire left_32_read_write_en;
  wire left_32_read_clk;
  wire [31:0] left_32_read_out;
  wire left_32_read_done;
  wire [31:0] top_32_read_in;
  wire top_32_read_write_en;
  wire top_32_read_clk;
  wire [31:0] top_32_read_out;
  wire top_32_read_done;
  wire [31:0] pe_32_top;
  wire [31:0] pe_32_left;
  wire pe_32_go;
  wire pe_32_clk;
  wire [31:0] pe_32_down;
  wire [31:0] pe_32_right;
  wire [31:0] pe_32_out;
  wire pe_32_done;
  wire [31:0] down_31_write_in;
  wire down_31_write_write_en;
  wire down_31_write_clk;
  wire [31:0] down_31_write_out;
  wire down_31_write_done;
  wire [31:0] right_31_write_in;
  wire right_31_write_write_en;
  wire right_31_write_clk;
  wire [31:0] right_31_write_out;
  wire right_31_write_done;
  wire [31:0] left_31_read_in;
  wire left_31_read_write_en;
  wire left_31_read_clk;
  wire [31:0] left_31_read_out;
  wire left_31_read_done;
  wire [31:0] top_31_read_in;
  wire top_31_read_write_en;
  wire top_31_read_clk;
  wire [31:0] top_31_read_out;
  wire top_31_read_done;
  wire [31:0] pe_31_top;
  wire [31:0] pe_31_left;
  wire pe_31_go;
  wire pe_31_clk;
  wire [31:0] pe_31_down;
  wire [31:0] pe_31_right;
  wire [31:0] pe_31_out;
  wire pe_31_done;
  wire [31:0] down_30_write_in;
  wire down_30_write_write_en;
  wire down_30_write_clk;
  wire [31:0] down_30_write_out;
  wire down_30_write_done;
  wire [31:0] right_30_write_in;
  wire right_30_write_write_en;
  wire right_30_write_clk;
  wire [31:0] right_30_write_out;
  wire right_30_write_done;
  wire [31:0] left_30_read_in;
  wire left_30_read_write_en;
  wire left_30_read_clk;
  wire [31:0] left_30_read_out;
  wire left_30_read_done;
  wire [31:0] top_30_read_in;
  wire top_30_read_write_en;
  wire top_30_read_clk;
  wire [31:0] top_30_read_out;
  wire top_30_read_done;
  wire [31:0] pe_30_top;
  wire [31:0] pe_30_left;
  wire pe_30_go;
  wire pe_30_clk;
  wire [31:0] pe_30_down;
  wire [31:0] pe_30_right;
  wire [31:0] pe_30_out;
  wire pe_30_done;
  wire [31:0] down_25_write_in;
  wire down_25_write_write_en;
  wire down_25_write_clk;
  wire [31:0] down_25_write_out;
  wire down_25_write_done;
  wire [31:0] left_25_read_in;
  wire left_25_read_write_en;
  wire left_25_read_clk;
  wire [31:0] left_25_read_out;
  wire left_25_read_done;
  wire [31:0] top_25_read_in;
  wire top_25_read_write_en;
  wire top_25_read_clk;
  wire [31:0] top_25_read_out;
  wire top_25_read_done;
  wire [31:0] pe_25_top;
  wire [31:0] pe_25_left;
  wire pe_25_go;
  wire pe_25_clk;
  wire [31:0] pe_25_down;
  wire [31:0] pe_25_right;
  wire [31:0] pe_25_out;
  wire pe_25_done;
  wire [31:0] down_24_write_in;
  wire down_24_write_write_en;
  wire down_24_write_clk;
  wire [31:0] down_24_write_out;
  wire down_24_write_done;
  wire [31:0] right_24_write_in;
  wire right_24_write_write_en;
  wire right_24_write_clk;
  wire [31:0] right_24_write_out;
  wire right_24_write_done;
  wire [31:0] left_24_read_in;
  wire left_24_read_write_en;
  wire left_24_read_clk;
  wire [31:0] left_24_read_out;
  wire left_24_read_done;
  wire [31:0] top_24_read_in;
  wire top_24_read_write_en;
  wire top_24_read_clk;
  wire [31:0] top_24_read_out;
  wire top_24_read_done;
  wire [31:0] pe_24_top;
  wire [31:0] pe_24_left;
  wire pe_24_go;
  wire pe_24_clk;
  wire [31:0] pe_24_down;
  wire [31:0] pe_24_right;
  wire [31:0] pe_24_out;
  wire pe_24_done;
  wire [31:0] down_23_write_in;
  wire down_23_write_write_en;
  wire down_23_write_clk;
  wire [31:0] down_23_write_out;
  wire down_23_write_done;
  wire [31:0] right_23_write_in;
  wire right_23_write_write_en;
  wire right_23_write_clk;
  wire [31:0] right_23_write_out;
  wire right_23_write_done;
  wire [31:0] left_23_read_in;
  wire left_23_read_write_en;
  wire left_23_read_clk;
  wire [31:0] left_23_read_out;
  wire left_23_read_done;
  wire [31:0] top_23_read_in;
  wire top_23_read_write_en;
  wire top_23_read_clk;
  wire [31:0] top_23_read_out;
  wire top_23_read_done;
  wire [31:0] pe_23_top;
  wire [31:0] pe_23_left;
  wire pe_23_go;
  wire pe_23_clk;
  wire [31:0] pe_23_down;
  wire [31:0] pe_23_right;
  wire [31:0] pe_23_out;
  wire pe_23_done;
  wire [31:0] down_22_write_in;
  wire down_22_write_write_en;
  wire down_22_write_clk;
  wire [31:0] down_22_write_out;
  wire down_22_write_done;
  wire [31:0] right_22_write_in;
  wire right_22_write_write_en;
  wire right_22_write_clk;
  wire [31:0] right_22_write_out;
  wire right_22_write_done;
  wire [31:0] left_22_read_in;
  wire left_22_read_write_en;
  wire left_22_read_clk;
  wire [31:0] left_22_read_out;
  wire left_22_read_done;
  wire [31:0] top_22_read_in;
  wire top_22_read_write_en;
  wire top_22_read_clk;
  wire [31:0] top_22_read_out;
  wire top_22_read_done;
  wire [31:0] pe_22_top;
  wire [31:0] pe_22_left;
  wire pe_22_go;
  wire pe_22_clk;
  wire [31:0] pe_22_down;
  wire [31:0] pe_22_right;
  wire [31:0] pe_22_out;
  wire pe_22_done;
  wire [31:0] down_21_write_in;
  wire down_21_write_write_en;
  wire down_21_write_clk;
  wire [31:0] down_21_write_out;
  wire down_21_write_done;
  wire [31:0] right_21_write_in;
  wire right_21_write_write_en;
  wire right_21_write_clk;
  wire [31:0] right_21_write_out;
  wire right_21_write_done;
  wire [31:0] left_21_read_in;
  wire left_21_read_write_en;
  wire left_21_read_clk;
  wire [31:0] left_21_read_out;
  wire left_21_read_done;
  wire [31:0] top_21_read_in;
  wire top_21_read_write_en;
  wire top_21_read_clk;
  wire [31:0] top_21_read_out;
  wire top_21_read_done;
  wire [31:0] pe_21_top;
  wire [31:0] pe_21_left;
  wire pe_21_go;
  wire pe_21_clk;
  wire [31:0] pe_21_down;
  wire [31:0] pe_21_right;
  wire [31:0] pe_21_out;
  wire pe_21_done;
  wire [31:0] down_20_write_in;
  wire down_20_write_write_en;
  wire down_20_write_clk;
  wire [31:0] down_20_write_out;
  wire down_20_write_done;
  wire [31:0] right_20_write_in;
  wire right_20_write_write_en;
  wire right_20_write_clk;
  wire [31:0] right_20_write_out;
  wire right_20_write_done;
  wire [31:0] left_20_read_in;
  wire left_20_read_write_en;
  wire left_20_read_clk;
  wire [31:0] left_20_read_out;
  wire left_20_read_done;
  wire [31:0] top_20_read_in;
  wire top_20_read_write_en;
  wire top_20_read_clk;
  wire [31:0] top_20_read_out;
  wire top_20_read_done;
  wire [31:0] pe_20_top;
  wire [31:0] pe_20_left;
  wire pe_20_go;
  wire pe_20_clk;
  wire [31:0] pe_20_down;
  wire [31:0] pe_20_right;
  wire [31:0] pe_20_out;
  wire pe_20_done;
  wire [31:0] down_15_write_in;
  wire down_15_write_write_en;
  wire down_15_write_clk;
  wire [31:0] down_15_write_out;
  wire down_15_write_done;
  wire [31:0] left_15_read_in;
  wire left_15_read_write_en;
  wire left_15_read_clk;
  wire [31:0] left_15_read_out;
  wire left_15_read_done;
  wire [31:0] top_15_read_in;
  wire top_15_read_write_en;
  wire top_15_read_clk;
  wire [31:0] top_15_read_out;
  wire top_15_read_done;
  wire [31:0] pe_15_top;
  wire [31:0] pe_15_left;
  wire pe_15_go;
  wire pe_15_clk;
  wire [31:0] pe_15_down;
  wire [31:0] pe_15_right;
  wire [31:0] pe_15_out;
  wire pe_15_done;
  wire [31:0] down_14_write_in;
  wire down_14_write_write_en;
  wire down_14_write_clk;
  wire [31:0] down_14_write_out;
  wire down_14_write_done;
  wire [31:0] right_14_write_in;
  wire right_14_write_write_en;
  wire right_14_write_clk;
  wire [31:0] right_14_write_out;
  wire right_14_write_done;
  wire [31:0] left_14_read_in;
  wire left_14_read_write_en;
  wire left_14_read_clk;
  wire [31:0] left_14_read_out;
  wire left_14_read_done;
  wire [31:0] top_14_read_in;
  wire top_14_read_write_en;
  wire top_14_read_clk;
  wire [31:0] top_14_read_out;
  wire top_14_read_done;
  wire [31:0] pe_14_top;
  wire [31:0] pe_14_left;
  wire pe_14_go;
  wire pe_14_clk;
  wire [31:0] pe_14_down;
  wire [31:0] pe_14_right;
  wire [31:0] pe_14_out;
  wire pe_14_done;
  wire [31:0] down_13_write_in;
  wire down_13_write_write_en;
  wire down_13_write_clk;
  wire [31:0] down_13_write_out;
  wire down_13_write_done;
  wire [31:0] right_13_write_in;
  wire right_13_write_write_en;
  wire right_13_write_clk;
  wire [31:0] right_13_write_out;
  wire right_13_write_done;
  wire [31:0] left_13_read_in;
  wire left_13_read_write_en;
  wire left_13_read_clk;
  wire [31:0] left_13_read_out;
  wire left_13_read_done;
  wire [31:0] top_13_read_in;
  wire top_13_read_write_en;
  wire top_13_read_clk;
  wire [31:0] top_13_read_out;
  wire top_13_read_done;
  wire [31:0] pe_13_top;
  wire [31:0] pe_13_left;
  wire pe_13_go;
  wire pe_13_clk;
  wire [31:0] pe_13_down;
  wire [31:0] pe_13_right;
  wire [31:0] pe_13_out;
  wire pe_13_done;
  wire [31:0] down_12_write_in;
  wire down_12_write_write_en;
  wire down_12_write_clk;
  wire [31:0] down_12_write_out;
  wire down_12_write_done;
  wire [31:0] right_12_write_in;
  wire right_12_write_write_en;
  wire right_12_write_clk;
  wire [31:0] right_12_write_out;
  wire right_12_write_done;
  wire [31:0] left_12_read_in;
  wire left_12_read_write_en;
  wire left_12_read_clk;
  wire [31:0] left_12_read_out;
  wire left_12_read_done;
  wire [31:0] top_12_read_in;
  wire top_12_read_write_en;
  wire top_12_read_clk;
  wire [31:0] top_12_read_out;
  wire top_12_read_done;
  wire [31:0] pe_12_top;
  wire [31:0] pe_12_left;
  wire pe_12_go;
  wire pe_12_clk;
  wire [31:0] pe_12_down;
  wire [31:0] pe_12_right;
  wire [31:0] pe_12_out;
  wire pe_12_done;
  wire [31:0] down_11_write_in;
  wire down_11_write_write_en;
  wire down_11_write_clk;
  wire [31:0] down_11_write_out;
  wire down_11_write_done;
  wire [31:0] right_11_write_in;
  wire right_11_write_write_en;
  wire right_11_write_clk;
  wire [31:0] right_11_write_out;
  wire right_11_write_done;
  wire [31:0] left_11_read_in;
  wire left_11_read_write_en;
  wire left_11_read_clk;
  wire [31:0] left_11_read_out;
  wire left_11_read_done;
  wire [31:0] top_11_read_in;
  wire top_11_read_write_en;
  wire top_11_read_clk;
  wire [31:0] top_11_read_out;
  wire top_11_read_done;
  wire [31:0] pe_11_top;
  wire [31:0] pe_11_left;
  wire pe_11_go;
  wire pe_11_clk;
  wire [31:0] pe_11_down;
  wire [31:0] pe_11_right;
  wire [31:0] pe_11_out;
  wire pe_11_done;
  wire [31:0] down_10_write_in;
  wire down_10_write_write_en;
  wire down_10_write_clk;
  wire [31:0] down_10_write_out;
  wire down_10_write_done;
  wire [31:0] right_10_write_in;
  wire right_10_write_write_en;
  wire right_10_write_clk;
  wire [31:0] right_10_write_out;
  wire right_10_write_done;
  wire [31:0] left_10_read_in;
  wire left_10_read_write_en;
  wire left_10_read_clk;
  wire [31:0] left_10_read_out;
  wire left_10_read_done;
  wire [31:0] top_10_read_in;
  wire top_10_read_write_en;
  wire top_10_read_clk;
  wire [31:0] top_10_read_out;
  wire top_10_read_done;
  wire [31:0] pe_10_top;
  wire [31:0] pe_10_left;
  wire pe_10_go;
  wire pe_10_clk;
  wire [31:0] pe_10_down;
  wire [31:0] pe_10_right;
  wire [31:0] pe_10_out;
  wire pe_10_done;
  wire [31:0] down_05_write_in;
  wire down_05_write_write_en;
  wire down_05_write_clk;
  wire [31:0] down_05_write_out;
  wire down_05_write_done;
  wire [31:0] left_05_read_in;
  wire left_05_read_write_en;
  wire left_05_read_clk;
  wire [31:0] left_05_read_out;
  wire left_05_read_done;
  wire [31:0] top_05_read_in;
  wire top_05_read_write_en;
  wire top_05_read_clk;
  wire [31:0] top_05_read_out;
  wire top_05_read_done;
  wire [31:0] pe_05_top;
  wire [31:0] pe_05_left;
  wire pe_05_go;
  wire pe_05_clk;
  wire [31:0] pe_05_down;
  wire [31:0] pe_05_right;
  wire [31:0] pe_05_out;
  wire pe_05_done;
  wire [31:0] down_04_write_in;
  wire down_04_write_write_en;
  wire down_04_write_clk;
  wire [31:0] down_04_write_out;
  wire down_04_write_done;
  wire [31:0] right_04_write_in;
  wire right_04_write_write_en;
  wire right_04_write_clk;
  wire [31:0] right_04_write_out;
  wire right_04_write_done;
  wire [31:0] left_04_read_in;
  wire left_04_read_write_en;
  wire left_04_read_clk;
  wire [31:0] left_04_read_out;
  wire left_04_read_done;
  wire [31:0] top_04_read_in;
  wire top_04_read_write_en;
  wire top_04_read_clk;
  wire [31:0] top_04_read_out;
  wire top_04_read_done;
  wire [31:0] pe_04_top;
  wire [31:0] pe_04_left;
  wire pe_04_go;
  wire pe_04_clk;
  wire [31:0] pe_04_down;
  wire [31:0] pe_04_right;
  wire [31:0] pe_04_out;
  wire pe_04_done;
  wire [31:0] down_03_write_in;
  wire down_03_write_write_en;
  wire down_03_write_clk;
  wire [31:0] down_03_write_out;
  wire down_03_write_done;
  wire [31:0] right_03_write_in;
  wire right_03_write_write_en;
  wire right_03_write_clk;
  wire [31:0] right_03_write_out;
  wire right_03_write_done;
  wire [31:0] left_03_read_in;
  wire left_03_read_write_en;
  wire left_03_read_clk;
  wire [31:0] left_03_read_out;
  wire left_03_read_done;
  wire [31:0] top_03_read_in;
  wire top_03_read_write_en;
  wire top_03_read_clk;
  wire [31:0] top_03_read_out;
  wire top_03_read_done;
  wire [31:0] pe_03_top;
  wire [31:0] pe_03_left;
  wire pe_03_go;
  wire pe_03_clk;
  wire [31:0] pe_03_down;
  wire [31:0] pe_03_right;
  wire [31:0] pe_03_out;
  wire pe_03_done;
  wire [31:0] down_02_write_in;
  wire down_02_write_write_en;
  wire down_02_write_clk;
  wire [31:0] down_02_write_out;
  wire down_02_write_done;
  wire [31:0] right_02_write_in;
  wire right_02_write_write_en;
  wire right_02_write_clk;
  wire [31:0] right_02_write_out;
  wire right_02_write_done;
  wire [31:0] left_02_read_in;
  wire left_02_read_write_en;
  wire left_02_read_clk;
  wire [31:0] left_02_read_out;
  wire left_02_read_done;
  wire [31:0] top_02_read_in;
  wire top_02_read_write_en;
  wire top_02_read_clk;
  wire [31:0] top_02_read_out;
  wire top_02_read_done;
  wire [31:0] pe_02_top;
  wire [31:0] pe_02_left;
  wire pe_02_go;
  wire pe_02_clk;
  wire [31:0] pe_02_down;
  wire [31:0] pe_02_right;
  wire [31:0] pe_02_out;
  wire pe_02_done;
  wire [31:0] down_01_write_in;
  wire down_01_write_write_en;
  wire down_01_write_clk;
  wire [31:0] down_01_write_out;
  wire down_01_write_done;
  wire [31:0] right_01_write_in;
  wire right_01_write_write_en;
  wire right_01_write_clk;
  wire [31:0] right_01_write_out;
  wire right_01_write_done;
  wire [31:0] left_01_read_in;
  wire left_01_read_write_en;
  wire left_01_read_clk;
  wire [31:0] left_01_read_out;
  wire left_01_read_done;
  wire [31:0] top_01_read_in;
  wire top_01_read_write_en;
  wire top_01_read_clk;
  wire [31:0] top_01_read_out;
  wire top_01_read_done;
  wire [31:0] pe_01_top;
  wire [31:0] pe_01_left;
  wire pe_01_go;
  wire pe_01_clk;
  wire [31:0] pe_01_down;
  wire [31:0] pe_01_right;
  wire [31:0] pe_01_out;
  wire pe_01_done;
  wire [31:0] down_00_write_in;
  wire down_00_write_write_en;
  wire down_00_write_clk;
  wire [31:0] down_00_write_out;
  wire down_00_write_done;
  wire [31:0] right_00_write_in;
  wire right_00_write_write_en;
  wire right_00_write_clk;
  wire [31:0] right_00_write_out;
  wire right_00_write_done;
  wire [31:0] left_00_read_in;
  wire left_00_read_write_en;
  wire left_00_read_clk;
  wire [31:0] left_00_read_out;
  wire left_00_read_done;
  wire [31:0] top_00_read_in;
  wire top_00_read_write_en;
  wire top_00_read_clk;
  wire [31:0] top_00_read_out;
  wire top_00_read_done;
  wire [31:0] pe_00_top;
  wire [31:0] pe_00_left;
  wire pe_00_go;
  wire pe_00_clk;
  wire [31:0] pe_00_down;
  wire [31:0] pe_00_right;
  wire [31:0] pe_00_out;
  wire pe_00_done;
  wire [2:0] l5_addr0;
  wire [31:0] l5_write_data;
  wire l5_write_en;
  wire l5_clk;
  wire [31:0] l5_read_data;
  wire l5_done;
  wire [2:0] l5_add_left;
  wire [2:0] l5_add_right;
  wire [2:0] l5_add_out;
  wire [2:0] l5_idx_in;
  wire l5_idx_write_en;
  wire l5_idx_clk;
  wire [2:0] l5_idx_out;
  wire l5_idx_done;
  wire [2:0] l4_addr0;
  wire [31:0] l4_write_data;
  wire l4_write_en;
  wire l4_clk;
  wire [31:0] l4_read_data;
  wire l4_done;
  wire [2:0] l4_add_left;
  wire [2:0] l4_add_right;
  wire [2:0] l4_add_out;
  wire [2:0] l4_idx_in;
  wire l4_idx_write_en;
  wire l4_idx_clk;
  wire [2:0] l4_idx_out;
  wire l4_idx_done;
  wire [2:0] l3_addr0;
  wire [31:0] l3_write_data;
  wire l3_write_en;
  wire l3_clk;
  wire [31:0] l3_read_data;
  wire l3_done;
  wire [2:0] l3_add_left;
  wire [2:0] l3_add_right;
  wire [2:0] l3_add_out;
  wire [2:0] l3_idx_in;
  wire l3_idx_write_en;
  wire l3_idx_clk;
  wire [2:0] l3_idx_out;
  wire l3_idx_done;
  wire [2:0] l2_addr0;
  wire [31:0] l2_write_data;
  wire l2_write_en;
  wire l2_clk;
  wire [31:0] l2_read_data;
  wire l2_done;
  wire [2:0] l2_add_left;
  wire [2:0] l2_add_right;
  wire [2:0] l2_add_out;
  wire [2:0] l2_idx_in;
  wire l2_idx_write_en;
  wire l2_idx_clk;
  wire [2:0] l2_idx_out;
  wire l2_idx_done;
  wire [2:0] l1_addr0;
  wire [31:0] l1_write_data;
  wire l1_write_en;
  wire l1_clk;
  wire [31:0] l1_read_data;
  wire l1_done;
  wire [2:0] l1_add_left;
  wire [2:0] l1_add_right;
  wire [2:0] l1_add_out;
  wire [2:0] l1_idx_in;
  wire l1_idx_write_en;
  wire l1_idx_clk;
  wire [2:0] l1_idx_out;
  wire l1_idx_done;
  wire [2:0] l0_addr0;
  wire [31:0] l0_write_data;
  wire l0_write_en;
  wire l0_clk;
  wire [31:0] l0_read_data;
  wire l0_done;
  wire [2:0] l0_add_left;
  wire [2:0] l0_add_right;
  wire [2:0] l0_add_out;
  wire [2:0] l0_idx_in;
  wire l0_idx_write_en;
  wire l0_idx_clk;
  wire [2:0] l0_idx_out;
  wire l0_idx_done;
  wire [2:0] t5_addr0;
  wire [31:0] t5_write_data;
  wire t5_write_en;
  wire t5_clk;
  wire [31:0] t5_read_data;
  wire t5_done;
  wire [2:0] t5_add_left;
  wire [2:0] t5_add_right;
  wire [2:0] t5_add_out;
  wire [2:0] t5_idx_in;
  wire t5_idx_write_en;
  wire t5_idx_clk;
  wire [2:0] t5_idx_out;
  wire t5_idx_done;
  wire [2:0] t4_addr0;
  wire [31:0] t4_write_data;
  wire t4_write_en;
  wire t4_clk;
  wire [31:0] t4_read_data;
  wire t4_done;
  wire [2:0] t4_add_left;
  wire [2:0] t4_add_right;
  wire [2:0] t4_add_out;
  wire [2:0] t4_idx_in;
  wire t4_idx_write_en;
  wire t4_idx_clk;
  wire [2:0] t4_idx_out;
  wire t4_idx_done;
  wire [2:0] t3_addr0;
  wire [31:0] t3_write_data;
  wire t3_write_en;
  wire t3_clk;
  wire [31:0] t3_read_data;
  wire t3_done;
  wire [2:0] t3_add_left;
  wire [2:0] t3_add_right;
  wire [2:0] t3_add_out;
  wire [2:0] t3_idx_in;
  wire t3_idx_write_en;
  wire t3_idx_clk;
  wire [2:0] t3_idx_out;
  wire t3_idx_done;
  wire [2:0] t2_addr0;
  wire [31:0] t2_write_data;
  wire t2_write_en;
  wire t2_clk;
  wire [31:0] t2_read_data;
  wire t2_done;
  wire [2:0] t2_add_left;
  wire [2:0] t2_add_right;
  wire [2:0] t2_add_out;
  wire [2:0] t2_idx_in;
  wire t2_idx_write_en;
  wire t2_idx_clk;
  wire [2:0] t2_idx_out;
  wire t2_idx_done;
  wire [2:0] t1_addr0;
  wire [31:0] t1_write_data;
  wire t1_write_en;
  wire t1_clk;
  wire [31:0] t1_read_data;
  wire t1_done;
  wire [2:0] t1_add_left;
  wire [2:0] t1_add_right;
  wire [2:0] t1_add_out;
  wire [2:0] t1_idx_in;
  wire t1_idx_write_en;
  wire t1_idx_clk;
  wire [2:0] t1_idx_out;
  wire t1_idx_done;
  wire [2:0] t0_addr0;
  wire [31:0] t0_write_data;
  wire t0_write_en;
  wire t0_clk;
  wire [31:0] t0_read_data;
  wire t0_done;
  wire [2:0] t0_add_left;
  wire [2:0] t0_add_right;
  wire [2:0] t0_add_out;
  wire [2:0] t0_idx_in;
  wire t0_idx_write_en;
  wire t0_idx_clk;
  wire [2:0] t0_idx_out;
  wire t0_idx_done;
  wire par_reset0_in;
  wire par_reset0_write_en;
  wire par_reset0_clk;
  wire par_reset0_out;
  wire par_reset0_done;
  wire par_done_reg0_in;
  wire par_done_reg0_write_en;
  wire par_done_reg0_clk;
  wire par_done_reg0_out;
  wire par_done_reg0_done;
  wire par_done_reg1_in;
  wire par_done_reg1_write_en;
  wire par_done_reg1_clk;
  wire par_done_reg1_out;
  wire par_done_reg1_done;
  wire par_done_reg2_in;
  wire par_done_reg2_write_en;
  wire par_done_reg2_clk;
  wire par_done_reg2_out;
  wire par_done_reg2_done;
  wire par_done_reg3_in;
  wire par_done_reg3_write_en;
  wire par_done_reg3_clk;
  wire par_done_reg3_out;
  wire par_done_reg3_done;
  wire par_done_reg4_in;
  wire par_done_reg4_write_en;
  wire par_done_reg4_clk;
  wire par_done_reg4_out;
  wire par_done_reg4_done;
  wire par_done_reg5_in;
  wire par_done_reg5_write_en;
  wire par_done_reg5_clk;
  wire par_done_reg5_out;
  wire par_done_reg5_done;
  wire par_done_reg6_in;
  wire par_done_reg6_write_en;
  wire par_done_reg6_clk;
  wire par_done_reg6_out;
  wire par_done_reg6_done;
  wire par_done_reg7_in;
  wire par_done_reg7_write_en;
  wire par_done_reg7_clk;
  wire par_done_reg7_out;
  wire par_done_reg7_done;
  wire par_done_reg8_in;
  wire par_done_reg8_write_en;
  wire par_done_reg8_clk;
  wire par_done_reg8_out;
  wire par_done_reg8_done;
  wire par_done_reg9_in;
  wire par_done_reg9_write_en;
  wire par_done_reg9_clk;
  wire par_done_reg9_out;
  wire par_done_reg9_done;
  wire par_done_reg10_in;
  wire par_done_reg10_write_en;
  wire par_done_reg10_clk;
  wire par_done_reg10_out;
  wire par_done_reg10_done;
  wire par_done_reg11_in;
  wire par_done_reg11_write_en;
  wire par_done_reg11_clk;
  wire par_done_reg11_out;
  wire par_done_reg11_done;
  wire par_reset1_in;
  wire par_reset1_write_en;
  wire par_reset1_clk;
  wire par_reset1_out;
  wire par_reset1_done;
  wire par_done_reg12_in;
  wire par_done_reg12_write_en;
  wire par_done_reg12_clk;
  wire par_done_reg12_out;
  wire par_done_reg12_done;
  wire par_done_reg13_in;
  wire par_done_reg13_write_en;
  wire par_done_reg13_clk;
  wire par_done_reg13_out;
  wire par_done_reg13_done;
  wire par_reset2_in;
  wire par_reset2_write_en;
  wire par_reset2_clk;
  wire par_reset2_out;
  wire par_reset2_done;
  wire par_done_reg14_in;
  wire par_done_reg14_write_en;
  wire par_done_reg14_clk;
  wire par_done_reg14_out;
  wire par_done_reg14_done;
  wire par_done_reg15_in;
  wire par_done_reg15_write_en;
  wire par_done_reg15_clk;
  wire par_done_reg15_out;
  wire par_done_reg15_done;
  wire par_reset3_in;
  wire par_reset3_write_en;
  wire par_reset3_clk;
  wire par_reset3_out;
  wire par_reset3_done;
  wire par_done_reg16_in;
  wire par_done_reg16_write_en;
  wire par_done_reg16_clk;
  wire par_done_reg16_out;
  wire par_done_reg16_done;
  wire par_done_reg17_in;
  wire par_done_reg17_write_en;
  wire par_done_reg17_clk;
  wire par_done_reg17_out;
  wire par_done_reg17_done;
  wire par_done_reg18_in;
  wire par_done_reg18_write_en;
  wire par_done_reg18_clk;
  wire par_done_reg18_out;
  wire par_done_reg18_done;
  wire par_done_reg19_in;
  wire par_done_reg19_write_en;
  wire par_done_reg19_clk;
  wire par_done_reg19_out;
  wire par_done_reg19_done;
  wire par_done_reg20_in;
  wire par_done_reg20_write_en;
  wire par_done_reg20_clk;
  wire par_done_reg20_out;
  wire par_done_reg20_done;
  wire par_reset4_in;
  wire par_reset4_write_en;
  wire par_reset4_clk;
  wire par_reset4_out;
  wire par_reset4_done;
  wire par_done_reg21_in;
  wire par_done_reg21_write_en;
  wire par_done_reg21_clk;
  wire par_done_reg21_out;
  wire par_done_reg21_done;
  wire par_done_reg22_in;
  wire par_done_reg22_write_en;
  wire par_done_reg22_clk;
  wire par_done_reg22_out;
  wire par_done_reg22_done;
  wire par_done_reg23_in;
  wire par_done_reg23_write_en;
  wire par_done_reg23_clk;
  wire par_done_reg23_out;
  wire par_done_reg23_done;
  wire par_done_reg24_in;
  wire par_done_reg24_write_en;
  wire par_done_reg24_clk;
  wire par_done_reg24_out;
  wire par_done_reg24_done;
  wire par_done_reg25_in;
  wire par_done_reg25_write_en;
  wire par_done_reg25_clk;
  wire par_done_reg25_out;
  wire par_done_reg25_done;
  wire par_done_reg26_in;
  wire par_done_reg26_write_en;
  wire par_done_reg26_clk;
  wire par_done_reg26_out;
  wire par_done_reg26_done;
  wire par_reset5_in;
  wire par_reset5_write_en;
  wire par_reset5_clk;
  wire par_reset5_out;
  wire par_reset5_done;
  wire par_done_reg27_in;
  wire par_done_reg27_write_en;
  wire par_done_reg27_clk;
  wire par_done_reg27_out;
  wire par_done_reg27_done;
  wire par_done_reg28_in;
  wire par_done_reg28_write_en;
  wire par_done_reg28_clk;
  wire par_done_reg28_out;
  wire par_done_reg28_done;
  wire par_done_reg29_in;
  wire par_done_reg29_write_en;
  wire par_done_reg29_clk;
  wire par_done_reg29_out;
  wire par_done_reg29_done;
  wire par_done_reg30_in;
  wire par_done_reg30_write_en;
  wire par_done_reg30_clk;
  wire par_done_reg30_out;
  wire par_done_reg30_done;
  wire par_done_reg31_in;
  wire par_done_reg31_write_en;
  wire par_done_reg31_clk;
  wire par_done_reg31_out;
  wire par_done_reg31_done;
  wire par_done_reg32_in;
  wire par_done_reg32_write_en;
  wire par_done_reg32_clk;
  wire par_done_reg32_out;
  wire par_done_reg32_done;
  wire par_done_reg33_in;
  wire par_done_reg33_write_en;
  wire par_done_reg33_clk;
  wire par_done_reg33_out;
  wire par_done_reg33_done;
  wire par_done_reg34_in;
  wire par_done_reg34_write_en;
  wire par_done_reg34_clk;
  wire par_done_reg34_out;
  wire par_done_reg34_done;
  wire par_done_reg35_in;
  wire par_done_reg35_write_en;
  wire par_done_reg35_clk;
  wire par_done_reg35_out;
  wire par_done_reg35_done;
  wire par_reset6_in;
  wire par_reset6_write_en;
  wire par_reset6_clk;
  wire par_reset6_out;
  wire par_reset6_done;
  wire par_done_reg36_in;
  wire par_done_reg36_write_en;
  wire par_done_reg36_clk;
  wire par_done_reg36_out;
  wire par_done_reg36_done;
  wire par_done_reg37_in;
  wire par_done_reg37_write_en;
  wire par_done_reg37_clk;
  wire par_done_reg37_out;
  wire par_done_reg37_done;
  wire par_done_reg38_in;
  wire par_done_reg38_write_en;
  wire par_done_reg38_clk;
  wire par_done_reg38_out;
  wire par_done_reg38_done;
  wire par_done_reg39_in;
  wire par_done_reg39_write_en;
  wire par_done_reg39_clk;
  wire par_done_reg39_out;
  wire par_done_reg39_done;
  wire par_done_reg40_in;
  wire par_done_reg40_write_en;
  wire par_done_reg40_clk;
  wire par_done_reg40_out;
  wire par_done_reg40_done;
  wire par_done_reg41_in;
  wire par_done_reg41_write_en;
  wire par_done_reg41_clk;
  wire par_done_reg41_out;
  wire par_done_reg41_done;
  wire par_done_reg42_in;
  wire par_done_reg42_write_en;
  wire par_done_reg42_clk;
  wire par_done_reg42_out;
  wire par_done_reg42_done;
  wire par_done_reg43_in;
  wire par_done_reg43_write_en;
  wire par_done_reg43_clk;
  wire par_done_reg43_out;
  wire par_done_reg43_done;
  wire par_done_reg44_in;
  wire par_done_reg44_write_en;
  wire par_done_reg44_clk;
  wire par_done_reg44_out;
  wire par_done_reg44_done;
  wire par_done_reg45_in;
  wire par_done_reg45_write_en;
  wire par_done_reg45_clk;
  wire par_done_reg45_out;
  wire par_done_reg45_done;
  wire par_done_reg46_in;
  wire par_done_reg46_write_en;
  wire par_done_reg46_clk;
  wire par_done_reg46_out;
  wire par_done_reg46_done;
  wire par_done_reg47_in;
  wire par_done_reg47_write_en;
  wire par_done_reg47_clk;
  wire par_done_reg47_out;
  wire par_done_reg47_done;
  wire par_reset7_in;
  wire par_reset7_write_en;
  wire par_reset7_clk;
  wire par_reset7_out;
  wire par_reset7_done;
  wire par_done_reg48_in;
  wire par_done_reg48_write_en;
  wire par_done_reg48_clk;
  wire par_done_reg48_out;
  wire par_done_reg48_done;
  wire par_done_reg49_in;
  wire par_done_reg49_write_en;
  wire par_done_reg49_clk;
  wire par_done_reg49_out;
  wire par_done_reg49_done;
  wire par_done_reg50_in;
  wire par_done_reg50_write_en;
  wire par_done_reg50_clk;
  wire par_done_reg50_out;
  wire par_done_reg50_done;
  wire par_done_reg51_in;
  wire par_done_reg51_write_en;
  wire par_done_reg51_clk;
  wire par_done_reg51_out;
  wire par_done_reg51_done;
  wire par_done_reg52_in;
  wire par_done_reg52_write_en;
  wire par_done_reg52_clk;
  wire par_done_reg52_out;
  wire par_done_reg52_done;
  wire par_done_reg53_in;
  wire par_done_reg53_write_en;
  wire par_done_reg53_clk;
  wire par_done_reg53_out;
  wire par_done_reg53_done;
  wire par_done_reg54_in;
  wire par_done_reg54_write_en;
  wire par_done_reg54_clk;
  wire par_done_reg54_out;
  wire par_done_reg54_done;
  wire par_done_reg55_in;
  wire par_done_reg55_write_en;
  wire par_done_reg55_clk;
  wire par_done_reg55_out;
  wire par_done_reg55_done;
  wire par_done_reg56_in;
  wire par_done_reg56_write_en;
  wire par_done_reg56_clk;
  wire par_done_reg56_out;
  wire par_done_reg56_done;
  wire par_done_reg57_in;
  wire par_done_reg57_write_en;
  wire par_done_reg57_clk;
  wire par_done_reg57_out;
  wire par_done_reg57_done;
  wire par_done_reg58_in;
  wire par_done_reg58_write_en;
  wire par_done_reg58_clk;
  wire par_done_reg58_out;
  wire par_done_reg58_done;
  wire par_done_reg59_in;
  wire par_done_reg59_write_en;
  wire par_done_reg59_clk;
  wire par_done_reg59_out;
  wire par_done_reg59_done;
  wire par_done_reg60_in;
  wire par_done_reg60_write_en;
  wire par_done_reg60_clk;
  wire par_done_reg60_out;
  wire par_done_reg60_done;
  wire par_done_reg61_in;
  wire par_done_reg61_write_en;
  wire par_done_reg61_clk;
  wire par_done_reg61_out;
  wire par_done_reg61_done;
  wire par_reset8_in;
  wire par_reset8_write_en;
  wire par_reset8_clk;
  wire par_reset8_out;
  wire par_reset8_done;
  wire par_done_reg62_in;
  wire par_done_reg62_write_en;
  wire par_done_reg62_clk;
  wire par_done_reg62_out;
  wire par_done_reg62_done;
  wire par_done_reg63_in;
  wire par_done_reg63_write_en;
  wire par_done_reg63_clk;
  wire par_done_reg63_out;
  wire par_done_reg63_done;
  wire par_done_reg64_in;
  wire par_done_reg64_write_en;
  wire par_done_reg64_clk;
  wire par_done_reg64_out;
  wire par_done_reg64_done;
  wire par_done_reg65_in;
  wire par_done_reg65_write_en;
  wire par_done_reg65_clk;
  wire par_done_reg65_out;
  wire par_done_reg65_done;
  wire par_done_reg66_in;
  wire par_done_reg66_write_en;
  wire par_done_reg66_clk;
  wire par_done_reg66_out;
  wire par_done_reg66_done;
  wire par_done_reg67_in;
  wire par_done_reg67_write_en;
  wire par_done_reg67_clk;
  wire par_done_reg67_out;
  wire par_done_reg67_done;
  wire par_done_reg68_in;
  wire par_done_reg68_write_en;
  wire par_done_reg68_clk;
  wire par_done_reg68_out;
  wire par_done_reg68_done;
  wire par_done_reg69_in;
  wire par_done_reg69_write_en;
  wire par_done_reg69_clk;
  wire par_done_reg69_out;
  wire par_done_reg69_done;
  wire par_done_reg70_in;
  wire par_done_reg70_write_en;
  wire par_done_reg70_clk;
  wire par_done_reg70_out;
  wire par_done_reg70_done;
  wire par_done_reg71_in;
  wire par_done_reg71_write_en;
  wire par_done_reg71_clk;
  wire par_done_reg71_out;
  wire par_done_reg71_done;
  wire par_done_reg72_in;
  wire par_done_reg72_write_en;
  wire par_done_reg72_clk;
  wire par_done_reg72_out;
  wire par_done_reg72_done;
  wire par_done_reg73_in;
  wire par_done_reg73_write_en;
  wire par_done_reg73_clk;
  wire par_done_reg73_out;
  wire par_done_reg73_done;
  wire par_done_reg74_in;
  wire par_done_reg74_write_en;
  wire par_done_reg74_clk;
  wire par_done_reg74_out;
  wire par_done_reg74_done;
  wire par_done_reg75_in;
  wire par_done_reg75_write_en;
  wire par_done_reg75_clk;
  wire par_done_reg75_out;
  wire par_done_reg75_done;
  wire par_done_reg76_in;
  wire par_done_reg76_write_en;
  wire par_done_reg76_clk;
  wire par_done_reg76_out;
  wire par_done_reg76_done;
  wire par_done_reg77_in;
  wire par_done_reg77_write_en;
  wire par_done_reg77_clk;
  wire par_done_reg77_out;
  wire par_done_reg77_done;
  wire par_done_reg78_in;
  wire par_done_reg78_write_en;
  wire par_done_reg78_clk;
  wire par_done_reg78_out;
  wire par_done_reg78_done;
  wire par_done_reg79_in;
  wire par_done_reg79_write_en;
  wire par_done_reg79_clk;
  wire par_done_reg79_out;
  wire par_done_reg79_done;
  wire par_done_reg80_in;
  wire par_done_reg80_write_en;
  wire par_done_reg80_clk;
  wire par_done_reg80_out;
  wire par_done_reg80_done;
  wire par_done_reg81_in;
  wire par_done_reg81_write_en;
  wire par_done_reg81_clk;
  wire par_done_reg81_out;
  wire par_done_reg81_done;
  wire par_reset9_in;
  wire par_reset9_write_en;
  wire par_reset9_clk;
  wire par_reset9_out;
  wire par_reset9_done;
  wire par_done_reg82_in;
  wire par_done_reg82_write_en;
  wire par_done_reg82_clk;
  wire par_done_reg82_out;
  wire par_done_reg82_done;
  wire par_done_reg83_in;
  wire par_done_reg83_write_en;
  wire par_done_reg83_clk;
  wire par_done_reg83_out;
  wire par_done_reg83_done;
  wire par_done_reg84_in;
  wire par_done_reg84_write_en;
  wire par_done_reg84_clk;
  wire par_done_reg84_out;
  wire par_done_reg84_done;
  wire par_done_reg85_in;
  wire par_done_reg85_write_en;
  wire par_done_reg85_clk;
  wire par_done_reg85_out;
  wire par_done_reg85_done;
  wire par_done_reg86_in;
  wire par_done_reg86_write_en;
  wire par_done_reg86_clk;
  wire par_done_reg86_out;
  wire par_done_reg86_done;
  wire par_done_reg87_in;
  wire par_done_reg87_write_en;
  wire par_done_reg87_clk;
  wire par_done_reg87_out;
  wire par_done_reg87_done;
  wire par_done_reg88_in;
  wire par_done_reg88_write_en;
  wire par_done_reg88_clk;
  wire par_done_reg88_out;
  wire par_done_reg88_done;
  wire par_done_reg89_in;
  wire par_done_reg89_write_en;
  wire par_done_reg89_clk;
  wire par_done_reg89_out;
  wire par_done_reg89_done;
  wire par_done_reg90_in;
  wire par_done_reg90_write_en;
  wire par_done_reg90_clk;
  wire par_done_reg90_out;
  wire par_done_reg90_done;
  wire par_done_reg91_in;
  wire par_done_reg91_write_en;
  wire par_done_reg91_clk;
  wire par_done_reg91_out;
  wire par_done_reg91_done;
  wire par_done_reg92_in;
  wire par_done_reg92_write_en;
  wire par_done_reg92_clk;
  wire par_done_reg92_out;
  wire par_done_reg92_done;
  wire par_done_reg93_in;
  wire par_done_reg93_write_en;
  wire par_done_reg93_clk;
  wire par_done_reg93_out;
  wire par_done_reg93_done;
  wire par_done_reg94_in;
  wire par_done_reg94_write_en;
  wire par_done_reg94_clk;
  wire par_done_reg94_out;
  wire par_done_reg94_done;
  wire par_done_reg95_in;
  wire par_done_reg95_write_en;
  wire par_done_reg95_clk;
  wire par_done_reg95_out;
  wire par_done_reg95_done;
  wire par_done_reg96_in;
  wire par_done_reg96_write_en;
  wire par_done_reg96_clk;
  wire par_done_reg96_out;
  wire par_done_reg96_done;
  wire par_done_reg97_in;
  wire par_done_reg97_write_en;
  wire par_done_reg97_clk;
  wire par_done_reg97_out;
  wire par_done_reg97_done;
  wire par_done_reg98_in;
  wire par_done_reg98_write_en;
  wire par_done_reg98_clk;
  wire par_done_reg98_out;
  wire par_done_reg98_done;
  wire par_done_reg99_in;
  wire par_done_reg99_write_en;
  wire par_done_reg99_clk;
  wire par_done_reg99_out;
  wire par_done_reg99_done;
  wire par_done_reg100_in;
  wire par_done_reg100_write_en;
  wire par_done_reg100_clk;
  wire par_done_reg100_out;
  wire par_done_reg100_done;
  wire par_done_reg101_in;
  wire par_done_reg101_write_en;
  wire par_done_reg101_clk;
  wire par_done_reg101_out;
  wire par_done_reg101_done;
  wire par_reset10_in;
  wire par_reset10_write_en;
  wire par_reset10_clk;
  wire par_reset10_out;
  wire par_reset10_done;
  wire par_done_reg102_in;
  wire par_done_reg102_write_en;
  wire par_done_reg102_clk;
  wire par_done_reg102_out;
  wire par_done_reg102_done;
  wire par_done_reg103_in;
  wire par_done_reg103_write_en;
  wire par_done_reg103_clk;
  wire par_done_reg103_out;
  wire par_done_reg103_done;
  wire par_done_reg104_in;
  wire par_done_reg104_write_en;
  wire par_done_reg104_clk;
  wire par_done_reg104_out;
  wire par_done_reg104_done;
  wire par_done_reg105_in;
  wire par_done_reg105_write_en;
  wire par_done_reg105_clk;
  wire par_done_reg105_out;
  wire par_done_reg105_done;
  wire par_done_reg106_in;
  wire par_done_reg106_write_en;
  wire par_done_reg106_clk;
  wire par_done_reg106_out;
  wire par_done_reg106_done;
  wire par_done_reg107_in;
  wire par_done_reg107_write_en;
  wire par_done_reg107_clk;
  wire par_done_reg107_out;
  wire par_done_reg107_done;
  wire par_done_reg108_in;
  wire par_done_reg108_write_en;
  wire par_done_reg108_clk;
  wire par_done_reg108_out;
  wire par_done_reg108_done;
  wire par_done_reg109_in;
  wire par_done_reg109_write_en;
  wire par_done_reg109_clk;
  wire par_done_reg109_out;
  wire par_done_reg109_done;
  wire par_done_reg110_in;
  wire par_done_reg110_write_en;
  wire par_done_reg110_clk;
  wire par_done_reg110_out;
  wire par_done_reg110_done;
  wire par_done_reg111_in;
  wire par_done_reg111_write_en;
  wire par_done_reg111_clk;
  wire par_done_reg111_out;
  wire par_done_reg111_done;
  wire par_done_reg112_in;
  wire par_done_reg112_write_en;
  wire par_done_reg112_clk;
  wire par_done_reg112_out;
  wire par_done_reg112_done;
  wire par_done_reg113_in;
  wire par_done_reg113_write_en;
  wire par_done_reg113_clk;
  wire par_done_reg113_out;
  wire par_done_reg113_done;
  wire par_done_reg114_in;
  wire par_done_reg114_write_en;
  wire par_done_reg114_clk;
  wire par_done_reg114_out;
  wire par_done_reg114_done;
  wire par_done_reg115_in;
  wire par_done_reg115_write_en;
  wire par_done_reg115_clk;
  wire par_done_reg115_out;
  wire par_done_reg115_done;
  wire par_done_reg116_in;
  wire par_done_reg116_write_en;
  wire par_done_reg116_clk;
  wire par_done_reg116_out;
  wire par_done_reg116_done;
  wire par_done_reg117_in;
  wire par_done_reg117_write_en;
  wire par_done_reg117_clk;
  wire par_done_reg117_out;
  wire par_done_reg117_done;
  wire par_done_reg118_in;
  wire par_done_reg118_write_en;
  wire par_done_reg118_clk;
  wire par_done_reg118_out;
  wire par_done_reg118_done;
  wire par_done_reg119_in;
  wire par_done_reg119_write_en;
  wire par_done_reg119_clk;
  wire par_done_reg119_out;
  wire par_done_reg119_done;
  wire par_done_reg120_in;
  wire par_done_reg120_write_en;
  wire par_done_reg120_clk;
  wire par_done_reg120_out;
  wire par_done_reg120_done;
  wire par_done_reg121_in;
  wire par_done_reg121_write_en;
  wire par_done_reg121_clk;
  wire par_done_reg121_out;
  wire par_done_reg121_done;
  wire par_done_reg122_in;
  wire par_done_reg122_write_en;
  wire par_done_reg122_clk;
  wire par_done_reg122_out;
  wire par_done_reg122_done;
  wire par_done_reg123_in;
  wire par_done_reg123_write_en;
  wire par_done_reg123_clk;
  wire par_done_reg123_out;
  wire par_done_reg123_done;
  wire par_done_reg124_in;
  wire par_done_reg124_write_en;
  wire par_done_reg124_clk;
  wire par_done_reg124_out;
  wire par_done_reg124_done;
  wire par_done_reg125_in;
  wire par_done_reg125_write_en;
  wire par_done_reg125_clk;
  wire par_done_reg125_out;
  wire par_done_reg125_done;
  wire par_done_reg126_in;
  wire par_done_reg126_write_en;
  wire par_done_reg126_clk;
  wire par_done_reg126_out;
  wire par_done_reg126_done;
  wire par_done_reg127_in;
  wire par_done_reg127_write_en;
  wire par_done_reg127_clk;
  wire par_done_reg127_out;
  wire par_done_reg127_done;
  wire par_done_reg128_in;
  wire par_done_reg128_write_en;
  wire par_done_reg128_clk;
  wire par_done_reg128_out;
  wire par_done_reg128_done;
  wire par_done_reg129_in;
  wire par_done_reg129_write_en;
  wire par_done_reg129_clk;
  wire par_done_reg129_out;
  wire par_done_reg129_done;
  wire par_done_reg130_in;
  wire par_done_reg130_write_en;
  wire par_done_reg130_clk;
  wire par_done_reg130_out;
  wire par_done_reg130_done;
  wire par_done_reg131_in;
  wire par_done_reg131_write_en;
  wire par_done_reg131_clk;
  wire par_done_reg131_out;
  wire par_done_reg131_done;
  wire par_reset11_in;
  wire par_reset11_write_en;
  wire par_reset11_clk;
  wire par_reset11_out;
  wire par_reset11_done;
  wire par_done_reg132_in;
  wire par_done_reg132_write_en;
  wire par_done_reg132_clk;
  wire par_done_reg132_out;
  wire par_done_reg132_done;
  wire par_done_reg133_in;
  wire par_done_reg133_write_en;
  wire par_done_reg133_clk;
  wire par_done_reg133_out;
  wire par_done_reg133_done;
  wire par_done_reg134_in;
  wire par_done_reg134_write_en;
  wire par_done_reg134_clk;
  wire par_done_reg134_out;
  wire par_done_reg134_done;
  wire par_done_reg135_in;
  wire par_done_reg135_write_en;
  wire par_done_reg135_clk;
  wire par_done_reg135_out;
  wire par_done_reg135_done;
  wire par_done_reg136_in;
  wire par_done_reg136_write_en;
  wire par_done_reg136_clk;
  wire par_done_reg136_out;
  wire par_done_reg136_done;
  wire par_done_reg137_in;
  wire par_done_reg137_write_en;
  wire par_done_reg137_clk;
  wire par_done_reg137_out;
  wire par_done_reg137_done;
  wire par_done_reg138_in;
  wire par_done_reg138_write_en;
  wire par_done_reg138_clk;
  wire par_done_reg138_out;
  wire par_done_reg138_done;
  wire par_done_reg139_in;
  wire par_done_reg139_write_en;
  wire par_done_reg139_clk;
  wire par_done_reg139_out;
  wire par_done_reg139_done;
  wire par_done_reg140_in;
  wire par_done_reg140_write_en;
  wire par_done_reg140_clk;
  wire par_done_reg140_out;
  wire par_done_reg140_done;
  wire par_done_reg141_in;
  wire par_done_reg141_write_en;
  wire par_done_reg141_clk;
  wire par_done_reg141_out;
  wire par_done_reg141_done;
  wire par_done_reg142_in;
  wire par_done_reg142_write_en;
  wire par_done_reg142_clk;
  wire par_done_reg142_out;
  wire par_done_reg142_done;
  wire par_done_reg143_in;
  wire par_done_reg143_write_en;
  wire par_done_reg143_clk;
  wire par_done_reg143_out;
  wire par_done_reg143_done;
  wire par_done_reg144_in;
  wire par_done_reg144_write_en;
  wire par_done_reg144_clk;
  wire par_done_reg144_out;
  wire par_done_reg144_done;
  wire par_done_reg145_in;
  wire par_done_reg145_write_en;
  wire par_done_reg145_clk;
  wire par_done_reg145_out;
  wire par_done_reg145_done;
  wire par_done_reg146_in;
  wire par_done_reg146_write_en;
  wire par_done_reg146_clk;
  wire par_done_reg146_out;
  wire par_done_reg146_done;
  wire par_done_reg147_in;
  wire par_done_reg147_write_en;
  wire par_done_reg147_clk;
  wire par_done_reg147_out;
  wire par_done_reg147_done;
  wire par_done_reg148_in;
  wire par_done_reg148_write_en;
  wire par_done_reg148_clk;
  wire par_done_reg148_out;
  wire par_done_reg148_done;
  wire par_done_reg149_in;
  wire par_done_reg149_write_en;
  wire par_done_reg149_clk;
  wire par_done_reg149_out;
  wire par_done_reg149_done;
  wire par_done_reg150_in;
  wire par_done_reg150_write_en;
  wire par_done_reg150_clk;
  wire par_done_reg150_out;
  wire par_done_reg150_done;
  wire par_done_reg151_in;
  wire par_done_reg151_write_en;
  wire par_done_reg151_clk;
  wire par_done_reg151_out;
  wire par_done_reg151_done;
  wire par_done_reg152_in;
  wire par_done_reg152_write_en;
  wire par_done_reg152_clk;
  wire par_done_reg152_out;
  wire par_done_reg152_done;
  wire par_done_reg153_in;
  wire par_done_reg153_write_en;
  wire par_done_reg153_clk;
  wire par_done_reg153_out;
  wire par_done_reg153_done;
  wire par_done_reg154_in;
  wire par_done_reg154_write_en;
  wire par_done_reg154_clk;
  wire par_done_reg154_out;
  wire par_done_reg154_done;
  wire par_done_reg155_in;
  wire par_done_reg155_write_en;
  wire par_done_reg155_clk;
  wire par_done_reg155_out;
  wire par_done_reg155_done;
  wire par_done_reg156_in;
  wire par_done_reg156_write_en;
  wire par_done_reg156_clk;
  wire par_done_reg156_out;
  wire par_done_reg156_done;
  wire par_done_reg157_in;
  wire par_done_reg157_write_en;
  wire par_done_reg157_clk;
  wire par_done_reg157_out;
  wire par_done_reg157_done;
  wire par_done_reg158_in;
  wire par_done_reg158_write_en;
  wire par_done_reg158_clk;
  wire par_done_reg158_out;
  wire par_done_reg158_done;
  wire par_reset12_in;
  wire par_reset12_write_en;
  wire par_reset12_clk;
  wire par_reset12_out;
  wire par_reset12_done;
  wire par_done_reg159_in;
  wire par_done_reg159_write_en;
  wire par_done_reg159_clk;
  wire par_done_reg159_out;
  wire par_done_reg159_done;
  wire par_done_reg160_in;
  wire par_done_reg160_write_en;
  wire par_done_reg160_clk;
  wire par_done_reg160_out;
  wire par_done_reg160_done;
  wire par_done_reg161_in;
  wire par_done_reg161_write_en;
  wire par_done_reg161_clk;
  wire par_done_reg161_out;
  wire par_done_reg161_done;
  wire par_done_reg162_in;
  wire par_done_reg162_write_en;
  wire par_done_reg162_clk;
  wire par_done_reg162_out;
  wire par_done_reg162_done;
  wire par_done_reg163_in;
  wire par_done_reg163_write_en;
  wire par_done_reg163_clk;
  wire par_done_reg163_out;
  wire par_done_reg163_done;
  wire par_done_reg164_in;
  wire par_done_reg164_write_en;
  wire par_done_reg164_clk;
  wire par_done_reg164_out;
  wire par_done_reg164_done;
  wire par_done_reg165_in;
  wire par_done_reg165_write_en;
  wire par_done_reg165_clk;
  wire par_done_reg165_out;
  wire par_done_reg165_done;
  wire par_done_reg166_in;
  wire par_done_reg166_write_en;
  wire par_done_reg166_clk;
  wire par_done_reg166_out;
  wire par_done_reg166_done;
  wire par_done_reg167_in;
  wire par_done_reg167_write_en;
  wire par_done_reg167_clk;
  wire par_done_reg167_out;
  wire par_done_reg167_done;
  wire par_done_reg168_in;
  wire par_done_reg168_write_en;
  wire par_done_reg168_clk;
  wire par_done_reg168_out;
  wire par_done_reg168_done;
  wire par_done_reg169_in;
  wire par_done_reg169_write_en;
  wire par_done_reg169_clk;
  wire par_done_reg169_out;
  wire par_done_reg169_done;
  wire par_done_reg170_in;
  wire par_done_reg170_write_en;
  wire par_done_reg170_clk;
  wire par_done_reg170_out;
  wire par_done_reg170_done;
  wire par_done_reg171_in;
  wire par_done_reg171_write_en;
  wire par_done_reg171_clk;
  wire par_done_reg171_out;
  wire par_done_reg171_done;
  wire par_done_reg172_in;
  wire par_done_reg172_write_en;
  wire par_done_reg172_clk;
  wire par_done_reg172_out;
  wire par_done_reg172_done;
  wire par_done_reg173_in;
  wire par_done_reg173_write_en;
  wire par_done_reg173_clk;
  wire par_done_reg173_out;
  wire par_done_reg173_done;
  wire par_done_reg174_in;
  wire par_done_reg174_write_en;
  wire par_done_reg174_clk;
  wire par_done_reg174_out;
  wire par_done_reg174_done;
  wire par_done_reg175_in;
  wire par_done_reg175_write_en;
  wire par_done_reg175_clk;
  wire par_done_reg175_out;
  wire par_done_reg175_done;
  wire par_done_reg176_in;
  wire par_done_reg176_write_en;
  wire par_done_reg176_clk;
  wire par_done_reg176_out;
  wire par_done_reg176_done;
  wire par_done_reg177_in;
  wire par_done_reg177_write_en;
  wire par_done_reg177_clk;
  wire par_done_reg177_out;
  wire par_done_reg177_done;
  wire par_done_reg178_in;
  wire par_done_reg178_write_en;
  wire par_done_reg178_clk;
  wire par_done_reg178_out;
  wire par_done_reg178_done;
  wire par_done_reg179_in;
  wire par_done_reg179_write_en;
  wire par_done_reg179_clk;
  wire par_done_reg179_out;
  wire par_done_reg179_done;
  wire par_done_reg180_in;
  wire par_done_reg180_write_en;
  wire par_done_reg180_clk;
  wire par_done_reg180_out;
  wire par_done_reg180_done;
  wire par_done_reg181_in;
  wire par_done_reg181_write_en;
  wire par_done_reg181_clk;
  wire par_done_reg181_out;
  wire par_done_reg181_done;
  wire par_done_reg182_in;
  wire par_done_reg182_write_en;
  wire par_done_reg182_clk;
  wire par_done_reg182_out;
  wire par_done_reg182_done;
  wire par_done_reg183_in;
  wire par_done_reg183_write_en;
  wire par_done_reg183_clk;
  wire par_done_reg183_out;
  wire par_done_reg183_done;
  wire par_done_reg184_in;
  wire par_done_reg184_write_en;
  wire par_done_reg184_clk;
  wire par_done_reg184_out;
  wire par_done_reg184_done;
  wire par_done_reg185_in;
  wire par_done_reg185_write_en;
  wire par_done_reg185_clk;
  wire par_done_reg185_out;
  wire par_done_reg185_done;
  wire par_done_reg186_in;
  wire par_done_reg186_write_en;
  wire par_done_reg186_clk;
  wire par_done_reg186_out;
  wire par_done_reg186_done;
  wire par_done_reg187_in;
  wire par_done_reg187_write_en;
  wire par_done_reg187_clk;
  wire par_done_reg187_out;
  wire par_done_reg187_done;
  wire par_done_reg188_in;
  wire par_done_reg188_write_en;
  wire par_done_reg188_clk;
  wire par_done_reg188_out;
  wire par_done_reg188_done;
  wire par_done_reg189_in;
  wire par_done_reg189_write_en;
  wire par_done_reg189_clk;
  wire par_done_reg189_out;
  wire par_done_reg189_done;
  wire par_done_reg190_in;
  wire par_done_reg190_write_en;
  wire par_done_reg190_clk;
  wire par_done_reg190_out;
  wire par_done_reg190_done;
  wire par_done_reg191_in;
  wire par_done_reg191_write_en;
  wire par_done_reg191_clk;
  wire par_done_reg191_out;
  wire par_done_reg191_done;
  wire par_done_reg192_in;
  wire par_done_reg192_write_en;
  wire par_done_reg192_clk;
  wire par_done_reg192_out;
  wire par_done_reg192_done;
  wire par_done_reg193_in;
  wire par_done_reg193_write_en;
  wire par_done_reg193_clk;
  wire par_done_reg193_out;
  wire par_done_reg193_done;
  wire par_done_reg194_in;
  wire par_done_reg194_write_en;
  wire par_done_reg194_clk;
  wire par_done_reg194_out;
  wire par_done_reg194_done;
  wire par_done_reg195_in;
  wire par_done_reg195_write_en;
  wire par_done_reg195_clk;
  wire par_done_reg195_out;
  wire par_done_reg195_done;
  wire par_done_reg196_in;
  wire par_done_reg196_write_en;
  wire par_done_reg196_clk;
  wire par_done_reg196_out;
  wire par_done_reg196_done;
  wire par_done_reg197_in;
  wire par_done_reg197_write_en;
  wire par_done_reg197_clk;
  wire par_done_reg197_out;
  wire par_done_reg197_done;
  wire par_done_reg198_in;
  wire par_done_reg198_write_en;
  wire par_done_reg198_clk;
  wire par_done_reg198_out;
  wire par_done_reg198_done;
  wire par_done_reg199_in;
  wire par_done_reg199_write_en;
  wire par_done_reg199_clk;
  wire par_done_reg199_out;
  wire par_done_reg199_done;
  wire par_done_reg200_in;
  wire par_done_reg200_write_en;
  wire par_done_reg200_clk;
  wire par_done_reg200_out;
  wire par_done_reg200_done;
  wire par_reset13_in;
  wire par_reset13_write_en;
  wire par_reset13_clk;
  wire par_reset13_out;
  wire par_reset13_done;
  wire par_done_reg201_in;
  wire par_done_reg201_write_en;
  wire par_done_reg201_clk;
  wire par_done_reg201_out;
  wire par_done_reg201_done;
  wire par_done_reg202_in;
  wire par_done_reg202_write_en;
  wire par_done_reg202_clk;
  wire par_done_reg202_out;
  wire par_done_reg202_done;
  wire par_done_reg203_in;
  wire par_done_reg203_write_en;
  wire par_done_reg203_clk;
  wire par_done_reg203_out;
  wire par_done_reg203_done;
  wire par_done_reg204_in;
  wire par_done_reg204_write_en;
  wire par_done_reg204_clk;
  wire par_done_reg204_out;
  wire par_done_reg204_done;
  wire par_done_reg205_in;
  wire par_done_reg205_write_en;
  wire par_done_reg205_clk;
  wire par_done_reg205_out;
  wire par_done_reg205_done;
  wire par_done_reg206_in;
  wire par_done_reg206_write_en;
  wire par_done_reg206_clk;
  wire par_done_reg206_out;
  wire par_done_reg206_done;
  wire par_done_reg207_in;
  wire par_done_reg207_write_en;
  wire par_done_reg207_clk;
  wire par_done_reg207_out;
  wire par_done_reg207_done;
  wire par_done_reg208_in;
  wire par_done_reg208_write_en;
  wire par_done_reg208_clk;
  wire par_done_reg208_out;
  wire par_done_reg208_done;
  wire par_done_reg209_in;
  wire par_done_reg209_write_en;
  wire par_done_reg209_clk;
  wire par_done_reg209_out;
  wire par_done_reg209_done;
  wire par_done_reg210_in;
  wire par_done_reg210_write_en;
  wire par_done_reg210_clk;
  wire par_done_reg210_out;
  wire par_done_reg210_done;
  wire par_done_reg211_in;
  wire par_done_reg211_write_en;
  wire par_done_reg211_clk;
  wire par_done_reg211_out;
  wire par_done_reg211_done;
  wire par_done_reg212_in;
  wire par_done_reg212_write_en;
  wire par_done_reg212_clk;
  wire par_done_reg212_out;
  wire par_done_reg212_done;
  wire par_done_reg213_in;
  wire par_done_reg213_write_en;
  wire par_done_reg213_clk;
  wire par_done_reg213_out;
  wire par_done_reg213_done;
  wire par_done_reg214_in;
  wire par_done_reg214_write_en;
  wire par_done_reg214_clk;
  wire par_done_reg214_out;
  wire par_done_reg214_done;
  wire par_done_reg215_in;
  wire par_done_reg215_write_en;
  wire par_done_reg215_clk;
  wire par_done_reg215_out;
  wire par_done_reg215_done;
  wire par_done_reg216_in;
  wire par_done_reg216_write_en;
  wire par_done_reg216_clk;
  wire par_done_reg216_out;
  wire par_done_reg216_done;
  wire par_done_reg217_in;
  wire par_done_reg217_write_en;
  wire par_done_reg217_clk;
  wire par_done_reg217_out;
  wire par_done_reg217_done;
  wire par_done_reg218_in;
  wire par_done_reg218_write_en;
  wire par_done_reg218_clk;
  wire par_done_reg218_out;
  wire par_done_reg218_done;
  wire par_done_reg219_in;
  wire par_done_reg219_write_en;
  wire par_done_reg219_clk;
  wire par_done_reg219_out;
  wire par_done_reg219_done;
  wire par_done_reg220_in;
  wire par_done_reg220_write_en;
  wire par_done_reg220_clk;
  wire par_done_reg220_out;
  wire par_done_reg220_done;
  wire par_done_reg221_in;
  wire par_done_reg221_write_en;
  wire par_done_reg221_clk;
  wire par_done_reg221_out;
  wire par_done_reg221_done;
  wire par_done_reg222_in;
  wire par_done_reg222_write_en;
  wire par_done_reg222_clk;
  wire par_done_reg222_out;
  wire par_done_reg222_done;
  wire par_done_reg223_in;
  wire par_done_reg223_write_en;
  wire par_done_reg223_clk;
  wire par_done_reg223_out;
  wire par_done_reg223_done;
  wire par_done_reg224_in;
  wire par_done_reg224_write_en;
  wire par_done_reg224_clk;
  wire par_done_reg224_out;
  wire par_done_reg224_done;
  wire par_done_reg225_in;
  wire par_done_reg225_write_en;
  wire par_done_reg225_clk;
  wire par_done_reg225_out;
  wire par_done_reg225_done;
  wire par_done_reg226_in;
  wire par_done_reg226_write_en;
  wire par_done_reg226_clk;
  wire par_done_reg226_out;
  wire par_done_reg226_done;
  wire par_done_reg227_in;
  wire par_done_reg227_write_en;
  wire par_done_reg227_clk;
  wire par_done_reg227_out;
  wire par_done_reg227_done;
  wire par_done_reg228_in;
  wire par_done_reg228_write_en;
  wire par_done_reg228_clk;
  wire par_done_reg228_out;
  wire par_done_reg228_done;
  wire par_done_reg229_in;
  wire par_done_reg229_write_en;
  wire par_done_reg229_clk;
  wire par_done_reg229_out;
  wire par_done_reg229_done;
  wire par_done_reg230_in;
  wire par_done_reg230_write_en;
  wire par_done_reg230_clk;
  wire par_done_reg230_out;
  wire par_done_reg230_done;
  wire par_done_reg231_in;
  wire par_done_reg231_write_en;
  wire par_done_reg231_clk;
  wire par_done_reg231_out;
  wire par_done_reg231_done;
  wire par_reset14_in;
  wire par_reset14_write_en;
  wire par_reset14_clk;
  wire par_reset14_out;
  wire par_reset14_done;
  wire par_done_reg232_in;
  wire par_done_reg232_write_en;
  wire par_done_reg232_clk;
  wire par_done_reg232_out;
  wire par_done_reg232_done;
  wire par_done_reg233_in;
  wire par_done_reg233_write_en;
  wire par_done_reg233_clk;
  wire par_done_reg233_out;
  wire par_done_reg233_done;
  wire par_done_reg234_in;
  wire par_done_reg234_write_en;
  wire par_done_reg234_clk;
  wire par_done_reg234_out;
  wire par_done_reg234_done;
  wire par_done_reg235_in;
  wire par_done_reg235_write_en;
  wire par_done_reg235_clk;
  wire par_done_reg235_out;
  wire par_done_reg235_done;
  wire par_done_reg236_in;
  wire par_done_reg236_write_en;
  wire par_done_reg236_clk;
  wire par_done_reg236_out;
  wire par_done_reg236_done;
  wire par_done_reg237_in;
  wire par_done_reg237_write_en;
  wire par_done_reg237_clk;
  wire par_done_reg237_out;
  wire par_done_reg237_done;
  wire par_done_reg238_in;
  wire par_done_reg238_write_en;
  wire par_done_reg238_clk;
  wire par_done_reg238_out;
  wire par_done_reg238_done;
  wire par_done_reg239_in;
  wire par_done_reg239_write_en;
  wire par_done_reg239_clk;
  wire par_done_reg239_out;
  wire par_done_reg239_done;
  wire par_done_reg240_in;
  wire par_done_reg240_write_en;
  wire par_done_reg240_clk;
  wire par_done_reg240_out;
  wire par_done_reg240_done;
  wire par_done_reg241_in;
  wire par_done_reg241_write_en;
  wire par_done_reg241_clk;
  wire par_done_reg241_out;
  wire par_done_reg241_done;
  wire par_done_reg242_in;
  wire par_done_reg242_write_en;
  wire par_done_reg242_clk;
  wire par_done_reg242_out;
  wire par_done_reg242_done;
  wire par_done_reg243_in;
  wire par_done_reg243_write_en;
  wire par_done_reg243_clk;
  wire par_done_reg243_out;
  wire par_done_reg243_done;
  wire par_done_reg244_in;
  wire par_done_reg244_write_en;
  wire par_done_reg244_clk;
  wire par_done_reg244_out;
  wire par_done_reg244_done;
  wire par_done_reg245_in;
  wire par_done_reg245_write_en;
  wire par_done_reg245_clk;
  wire par_done_reg245_out;
  wire par_done_reg245_done;
  wire par_done_reg246_in;
  wire par_done_reg246_write_en;
  wire par_done_reg246_clk;
  wire par_done_reg246_out;
  wire par_done_reg246_done;
  wire par_done_reg247_in;
  wire par_done_reg247_write_en;
  wire par_done_reg247_clk;
  wire par_done_reg247_out;
  wire par_done_reg247_done;
  wire par_done_reg248_in;
  wire par_done_reg248_write_en;
  wire par_done_reg248_clk;
  wire par_done_reg248_out;
  wire par_done_reg248_done;
  wire par_done_reg249_in;
  wire par_done_reg249_write_en;
  wire par_done_reg249_clk;
  wire par_done_reg249_out;
  wire par_done_reg249_done;
  wire par_done_reg250_in;
  wire par_done_reg250_write_en;
  wire par_done_reg250_clk;
  wire par_done_reg250_out;
  wire par_done_reg250_done;
  wire par_done_reg251_in;
  wire par_done_reg251_write_en;
  wire par_done_reg251_clk;
  wire par_done_reg251_out;
  wire par_done_reg251_done;
  wire par_done_reg252_in;
  wire par_done_reg252_write_en;
  wire par_done_reg252_clk;
  wire par_done_reg252_out;
  wire par_done_reg252_done;
  wire par_done_reg253_in;
  wire par_done_reg253_write_en;
  wire par_done_reg253_clk;
  wire par_done_reg253_out;
  wire par_done_reg253_done;
  wire par_done_reg254_in;
  wire par_done_reg254_write_en;
  wire par_done_reg254_clk;
  wire par_done_reg254_out;
  wire par_done_reg254_done;
  wire par_done_reg255_in;
  wire par_done_reg255_write_en;
  wire par_done_reg255_clk;
  wire par_done_reg255_out;
  wire par_done_reg255_done;
  wire par_done_reg256_in;
  wire par_done_reg256_write_en;
  wire par_done_reg256_clk;
  wire par_done_reg256_out;
  wire par_done_reg256_done;
  wire par_done_reg257_in;
  wire par_done_reg257_write_en;
  wire par_done_reg257_clk;
  wire par_done_reg257_out;
  wire par_done_reg257_done;
  wire par_done_reg258_in;
  wire par_done_reg258_write_en;
  wire par_done_reg258_clk;
  wire par_done_reg258_out;
  wire par_done_reg258_done;
  wire par_done_reg259_in;
  wire par_done_reg259_write_en;
  wire par_done_reg259_clk;
  wire par_done_reg259_out;
  wire par_done_reg259_done;
  wire par_done_reg260_in;
  wire par_done_reg260_write_en;
  wire par_done_reg260_clk;
  wire par_done_reg260_out;
  wire par_done_reg260_done;
  wire par_done_reg261_in;
  wire par_done_reg261_write_en;
  wire par_done_reg261_clk;
  wire par_done_reg261_out;
  wire par_done_reg261_done;
  wire par_done_reg262_in;
  wire par_done_reg262_write_en;
  wire par_done_reg262_clk;
  wire par_done_reg262_out;
  wire par_done_reg262_done;
  wire par_done_reg263_in;
  wire par_done_reg263_write_en;
  wire par_done_reg263_clk;
  wire par_done_reg263_out;
  wire par_done_reg263_done;
  wire par_done_reg264_in;
  wire par_done_reg264_write_en;
  wire par_done_reg264_clk;
  wire par_done_reg264_out;
  wire par_done_reg264_done;
  wire par_done_reg265_in;
  wire par_done_reg265_write_en;
  wire par_done_reg265_clk;
  wire par_done_reg265_out;
  wire par_done_reg265_done;
  wire par_done_reg266_in;
  wire par_done_reg266_write_en;
  wire par_done_reg266_clk;
  wire par_done_reg266_out;
  wire par_done_reg266_done;
  wire par_done_reg267_in;
  wire par_done_reg267_write_en;
  wire par_done_reg267_clk;
  wire par_done_reg267_out;
  wire par_done_reg267_done;
  wire par_done_reg268_in;
  wire par_done_reg268_write_en;
  wire par_done_reg268_clk;
  wire par_done_reg268_out;
  wire par_done_reg268_done;
  wire par_done_reg269_in;
  wire par_done_reg269_write_en;
  wire par_done_reg269_clk;
  wire par_done_reg269_out;
  wire par_done_reg269_done;
  wire par_done_reg270_in;
  wire par_done_reg270_write_en;
  wire par_done_reg270_clk;
  wire par_done_reg270_out;
  wire par_done_reg270_done;
  wire par_done_reg271_in;
  wire par_done_reg271_write_en;
  wire par_done_reg271_clk;
  wire par_done_reg271_out;
  wire par_done_reg271_done;
  wire par_done_reg272_in;
  wire par_done_reg272_write_en;
  wire par_done_reg272_clk;
  wire par_done_reg272_out;
  wire par_done_reg272_done;
  wire par_done_reg273_in;
  wire par_done_reg273_write_en;
  wire par_done_reg273_clk;
  wire par_done_reg273_out;
  wire par_done_reg273_done;
  wire par_done_reg274_in;
  wire par_done_reg274_write_en;
  wire par_done_reg274_clk;
  wire par_done_reg274_out;
  wire par_done_reg274_done;
  wire par_done_reg275_in;
  wire par_done_reg275_write_en;
  wire par_done_reg275_clk;
  wire par_done_reg275_out;
  wire par_done_reg275_done;
  wire par_done_reg276_in;
  wire par_done_reg276_write_en;
  wire par_done_reg276_clk;
  wire par_done_reg276_out;
  wire par_done_reg276_done;
  wire par_done_reg277_in;
  wire par_done_reg277_write_en;
  wire par_done_reg277_clk;
  wire par_done_reg277_out;
  wire par_done_reg277_done;
  wire par_done_reg278_in;
  wire par_done_reg278_write_en;
  wire par_done_reg278_clk;
  wire par_done_reg278_out;
  wire par_done_reg278_done;
  wire par_done_reg279_in;
  wire par_done_reg279_write_en;
  wire par_done_reg279_clk;
  wire par_done_reg279_out;
  wire par_done_reg279_done;
  wire par_done_reg280_in;
  wire par_done_reg280_write_en;
  wire par_done_reg280_clk;
  wire par_done_reg280_out;
  wire par_done_reg280_done;
  wire par_done_reg281_in;
  wire par_done_reg281_write_en;
  wire par_done_reg281_clk;
  wire par_done_reg281_out;
  wire par_done_reg281_done;
  wire par_reset15_in;
  wire par_reset15_write_en;
  wire par_reset15_clk;
  wire par_reset15_out;
  wire par_reset15_done;
  wire par_done_reg282_in;
  wire par_done_reg282_write_en;
  wire par_done_reg282_clk;
  wire par_done_reg282_out;
  wire par_done_reg282_done;
  wire par_done_reg283_in;
  wire par_done_reg283_write_en;
  wire par_done_reg283_clk;
  wire par_done_reg283_out;
  wire par_done_reg283_done;
  wire par_done_reg284_in;
  wire par_done_reg284_write_en;
  wire par_done_reg284_clk;
  wire par_done_reg284_out;
  wire par_done_reg284_done;
  wire par_done_reg285_in;
  wire par_done_reg285_write_en;
  wire par_done_reg285_clk;
  wire par_done_reg285_out;
  wire par_done_reg285_done;
  wire par_done_reg286_in;
  wire par_done_reg286_write_en;
  wire par_done_reg286_clk;
  wire par_done_reg286_out;
  wire par_done_reg286_done;
  wire par_done_reg287_in;
  wire par_done_reg287_write_en;
  wire par_done_reg287_clk;
  wire par_done_reg287_out;
  wire par_done_reg287_done;
  wire par_done_reg288_in;
  wire par_done_reg288_write_en;
  wire par_done_reg288_clk;
  wire par_done_reg288_out;
  wire par_done_reg288_done;
  wire par_done_reg289_in;
  wire par_done_reg289_write_en;
  wire par_done_reg289_clk;
  wire par_done_reg289_out;
  wire par_done_reg289_done;
  wire par_done_reg290_in;
  wire par_done_reg290_write_en;
  wire par_done_reg290_clk;
  wire par_done_reg290_out;
  wire par_done_reg290_done;
  wire par_done_reg291_in;
  wire par_done_reg291_write_en;
  wire par_done_reg291_clk;
  wire par_done_reg291_out;
  wire par_done_reg291_done;
  wire par_done_reg292_in;
  wire par_done_reg292_write_en;
  wire par_done_reg292_clk;
  wire par_done_reg292_out;
  wire par_done_reg292_done;
  wire par_done_reg293_in;
  wire par_done_reg293_write_en;
  wire par_done_reg293_clk;
  wire par_done_reg293_out;
  wire par_done_reg293_done;
  wire par_done_reg294_in;
  wire par_done_reg294_write_en;
  wire par_done_reg294_clk;
  wire par_done_reg294_out;
  wire par_done_reg294_done;
  wire par_done_reg295_in;
  wire par_done_reg295_write_en;
  wire par_done_reg295_clk;
  wire par_done_reg295_out;
  wire par_done_reg295_done;
  wire par_done_reg296_in;
  wire par_done_reg296_write_en;
  wire par_done_reg296_clk;
  wire par_done_reg296_out;
  wire par_done_reg296_done;
  wire par_done_reg297_in;
  wire par_done_reg297_write_en;
  wire par_done_reg297_clk;
  wire par_done_reg297_out;
  wire par_done_reg297_done;
  wire par_done_reg298_in;
  wire par_done_reg298_write_en;
  wire par_done_reg298_clk;
  wire par_done_reg298_out;
  wire par_done_reg298_done;
  wire par_done_reg299_in;
  wire par_done_reg299_write_en;
  wire par_done_reg299_clk;
  wire par_done_reg299_out;
  wire par_done_reg299_done;
  wire par_done_reg300_in;
  wire par_done_reg300_write_en;
  wire par_done_reg300_clk;
  wire par_done_reg300_out;
  wire par_done_reg300_done;
  wire par_done_reg301_in;
  wire par_done_reg301_write_en;
  wire par_done_reg301_clk;
  wire par_done_reg301_out;
  wire par_done_reg301_done;
  wire par_done_reg302_in;
  wire par_done_reg302_write_en;
  wire par_done_reg302_clk;
  wire par_done_reg302_out;
  wire par_done_reg302_done;
  wire par_done_reg303_in;
  wire par_done_reg303_write_en;
  wire par_done_reg303_clk;
  wire par_done_reg303_out;
  wire par_done_reg303_done;
  wire par_done_reg304_in;
  wire par_done_reg304_write_en;
  wire par_done_reg304_clk;
  wire par_done_reg304_out;
  wire par_done_reg304_done;
  wire par_done_reg305_in;
  wire par_done_reg305_write_en;
  wire par_done_reg305_clk;
  wire par_done_reg305_out;
  wire par_done_reg305_done;
  wire par_done_reg306_in;
  wire par_done_reg306_write_en;
  wire par_done_reg306_clk;
  wire par_done_reg306_out;
  wire par_done_reg306_done;
  wire par_done_reg307_in;
  wire par_done_reg307_write_en;
  wire par_done_reg307_clk;
  wire par_done_reg307_out;
  wire par_done_reg307_done;
  wire par_done_reg308_in;
  wire par_done_reg308_write_en;
  wire par_done_reg308_clk;
  wire par_done_reg308_out;
  wire par_done_reg308_done;
  wire par_done_reg309_in;
  wire par_done_reg309_write_en;
  wire par_done_reg309_clk;
  wire par_done_reg309_out;
  wire par_done_reg309_done;
  wire par_done_reg310_in;
  wire par_done_reg310_write_en;
  wire par_done_reg310_clk;
  wire par_done_reg310_out;
  wire par_done_reg310_done;
  wire par_done_reg311_in;
  wire par_done_reg311_write_en;
  wire par_done_reg311_clk;
  wire par_done_reg311_out;
  wire par_done_reg311_done;
  wire par_done_reg312_in;
  wire par_done_reg312_write_en;
  wire par_done_reg312_clk;
  wire par_done_reg312_out;
  wire par_done_reg312_done;
  wire par_done_reg313_in;
  wire par_done_reg313_write_en;
  wire par_done_reg313_clk;
  wire par_done_reg313_out;
  wire par_done_reg313_done;
  wire par_done_reg314_in;
  wire par_done_reg314_write_en;
  wire par_done_reg314_clk;
  wire par_done_reg314_out;
  wire par_done_reg314_done;
  wire par_reset16_in;
  wire par_reset16_write_en;
  wire par_reset16_clk;
  wire par_reset16_out;
  wire par_reset16_done;
  wire par_done_reg315_in;
  wire par_done_reg315_write_en;
  wire par_done_reg315_clk;
  wire par_done_reg315_out;
  wire par_done_reg315_done;
  wire par_done_reg316_in;
  wire par_done_reg316_write_en;
  wire par_done_reg316_clk;
  wire par_done_reg316_out;
  wire par_done_reg316_done;
  wire par_done_reg317_in;
  wire par_done_reg317_write_en;
  wire par_done_reg317_clk;
  wire par_done_reg317_out;
  wire par_done_reg317_done;
  wire par_done_reg318_in;
  wire par_done_reg318_write_en;
  wire par_done_reg318_clk;
  wire par_done_reg318_out;
  wire par_done_reg318_done;
  wire par_done_reg319_in;
  wire par_done_reg319_write_en;
  wire par_done_reg319_clk;
  wire par_done_reg319_out;
  wire par_done_reg319_done;
  wire par_done_reg320_in;
  wire par_done_reg320_write_en;
  wire par_done_reg320_clk;
  wire par_done_reg320_out;
  wire par_done_reg320_done;
  wire par_done_reg321_in;
  wire par_done_reg321_write_en;
  wire par_done_reg321_clk;
  wire par_done_reg321_out;
  wire par_done_reg321_done;
  wire par_done_reg322_in;
  wire par_done_reg322_write_en;
  wire par_done_reg322_clk;
  wire par_done_reg322_out;
  wire par_done_reg322_done;
  wire par_done_reg323_in;
  wire par_done_reg323_write_en;
  wire par_done_reg323_clk;
  wire par_done_reg323_out;
  wire par_done_reg323_done;
  wire par_done_reg324_in;
  wire par_done_reg324_write_en;
  wire par_done_reg324_clk;
  wire par_done_reg324_out;
  wire par_done_reg324_done;
  wire par_done_reg325_in;
  wire par_done_reg325_write_en;
  wire par_done_reg325_clk;
  wire par_done_reg325_out;
  wire par_done_reg325_done;
  wire par_done_reg326_in;
  wire par_done_reg326_write_en;
  wire par_done_reg326_clk;
  wire par_done_reg326_out;
  wire par_done_reg326_done;
  wire par_done_reg327_in;
  wire par_done_reg327_write_en;
  wire par_done_reg327_clk;
  wire par_done_reg327_out;
  wire par_done_reg327_done;
  wire par_done_reg328_in;
  wire par_done_reg328_write_en;
  wire par_done_reg328_clk;
  wire par_done_reg328_out;
  wire par_done_reg328_done;
  wire par_done_reg329_in;
  wire par_done_reg329_write_en;
  wire par_done_reg329_clk;
  wire par_done_reg329_out;
  wire par_done_reg329_done;
  wire par_done_reg330_in;
  wire par_done_reg330_write_en;
  wire par_done_reg330_clk;
  wire par_done_reg330_out;
  wire par_done_reg330_done;
  wire par_done_reg331_in;
  wire par_done_reg331_write_en;
  wire par_done_reg331_clk;
  wire par_done_reg331_out;
  wire par_done_reg331_done;
  wire par_done_reg332_in;
  wire par_done_reg332_write_en;
  wire par_done_reg332_clk;
  wire par_done_reg332_out;
  wire par_done_reg332_done;
  wire par_done_reg333_in;
  wire par_done_reg333_write_en;
  wire par_done_reg333_clk;
  wire par_done_reg333_out;
  wire par_done_reg333_done;
  wire par_done_reg334_in;
  wire par_done_reg334_write_en;
  wire par_done_reg334_clk;
  wire par_done_reg334_out;
  wire par_done_reg334_done;
  wire par_done_reg335_in;
  wire par_done_reg335_write_en;
  wire par_done_reg335_clk;
  wire par_done_reg335_out;
  wire par_done_reg335_done;
  wire par_done_reg336_in;
  wire par_done_reg336_write_en;
  wire par_done_reg336_clk;
  wire par_done_reg336_out;
  wire par_done_reg336_done;
  wire par_done_reg337_in;
  wire par_done_reg337_write_en;
  wire par_done_reg337_clk;
  wire par_done_reg337_out;
  wire par_done_reg337_done;
  wire par_done_reg338_in;
  wire par_done_reg338_write_en;
  wire par_done_reg338_clk;
  wire par_done_reg338_out;
  wire par_done_reg338_done;
  wire par_done_reg339_in;
  wire par_done_reg339_write_en;
  wire par_done_reg339_clk;
  wire par_done_reg339_out;
  wire par_done_reg339_done;
  wire par_done_reg340_in;
  wire par_done_reg340_write_en;
  wire par_done_reg340_clk;
  wire par_done_reg340_out;
  wire par_done_reg340_done;
  wire par_done_reg341_in;
  wire par_done_reg341_write_en;
  wire par_done_reg341_clk;
  wire par_done_reg341_out;
  wire par_done_reg341_done;
  wire par_done_reg342_in;
  wire par_done_reg342_write_en;
  wire par_done_reg342_clk;
  wire par_done_reg342_out;
  wire par_done_reg342_done;
  wire par_done_reg343_in;
  wire par_done_reg343_write_en;
  wire par_done_reg343_clk;
  wire par_done_reg343_out;
  wire par_done_reg343_done;
  wire par_done_reg344_in;
  wire par_done_reg344_write_en;
  wire par_done_reg344_clk;
  wire par_done_reg344_out;
  wire par_done_reg344_done;
  wire par_done_reg345_in;
  wire par_done_reg345_write_en;
  wire par_done_reg345_clk;
  wire par_done_reg345_out;
  wire par_done_reg345_done;
  wire par_done_reg346_in;
  wire par_done_reg346_write_en;
  wire par_done_reg346_clk;
  wire par_done_reg346_out;
  wire par_done_reg346_done;
  wire par_done_reg347_in;
  wire par_done_reg347_write_en;
  wire par_done_reg347_clk;
  wire par_done_reg347_out;
  wire par_done_reg347_done;
  wire par_done_reg348_in;
  wire par_done_reg348_write_en;
  wire par_done_reg348_clk;
  wire par_done_reg348_out;
  wire par_done_reg348_done;
  wire par_done_reg349_in;
  wire par_done_reg349_write_en;
  wire par_done_reg349_clk;
  wire par_done_reg349_out;
  wire par_done_reg349_done;
  wire par_done_reg350_in;
  wire par_done_reg350_write_en;
  wire par_done_reg350_clk;
  wire par_done_reg350_out;
  wire par_done_reg350_done;
  wire par_done_reg351_in;
  wire par_done_reg351_write_en;
  wire par_done_reg351_clk;
  wire par_done_reg351_out;
  wire par_done_reg351_done;
  wire par_done_reg352_in;
  wire par_done_reg352_write_en;
  wire par_done_reg352_clk;
  wire par_done_reg352_out;
  wire par_done_reg352_done;
  wire par_done_reg353_in;
  wire par_done_reg353_write_en;
  wire par_done_reg353_clk;
  wire par_done_reg353_out;
  wire par_done_reg353_done;
  wire par_done_reg354_in;
  wire par_done_reg354_write_en;
  wire par_done_reg354_clk;
  wire par_done_reg354_out;
  wire par_done_reg354_done;
  wire par_done_reg355_in;
  wire par_done_reg355_write_en;
  wire par_done_reg355_clk;
  wire par_done_reg355_out;
  wire par_done_reg355_done;
  wire par_done_reg356_in;
  wire par_done_reg356_write_en;
  wire par_done_reg356_clk;
  wire par_done_reg356_out;
  wire par_done_reg356_done;
  wire par_done_reg357_in;
  wire par_done_reg357_write_en;
  wire par_done_reg357_clk;
  wire par_done_reg357_out;
  wire par_done_reg357_done;
  wire par_done_reg358_in;
  wire par_done_reg358_write_en;
  wire par_done_reg358_clk;
  wire par_done_reg358_out;
  wire par_done_reg358_done;
  wire par_done_reg359_in;
  wire par_done_reg359_write_en;
  wire par_done_reg359_clk;
  wire par_done_reg359_out;
  wire par_done_reg359_done;
  wire par_done_reg360_in;
  wire par_done_reg360_write_en;
  wire par_done_reg360_clk;
  wire par_done_reg360_out;
  wire par_done_reg360_done;
  wire par_done_reg361_in;
  wire par_done_reg361_write_en;
  wire par_done_reg361_clk;
  wire par_done_reg361_out;
  wire par_done_reg361_done;
  wire par_done_reg362_in;
  wire par_done_reg362_write_en;
  wire par_done_reg362_clk;
  wire par_done_reg362_out;
  wire par_done_reg362_done;
  wire par_done_reg363_in;
  wire par_done_reg363_write_en;
  wire par_done_reg363_clk;
  wire par_done_reg363_out;
  wire par_done_reg363_done;
  wire par_done_reg364_in;
  wire par_done_reg364_write_en;
  wire par_done_reg364_clk;
  wire par_done_reg364_out;
  wire par_done_reg364_done;
  wire par_done_reg365_in;
  wire par_done_reg365_write_en;
  wire par_done_reg365_clk;
  wire par_done_reg365_out;
  wire par_done_reg365_done;
  wire par_done_reg366_in;
  wire par_done_reg366_write_en;
  wire par_done_reg366_clk;
  wire par_done_reg366_out;
  wire par_done_reg366_done;
  wire par_done_reg367_in;
  wire par_done_reg367_write_en;
  wire par_done_reg367_clk;
  wire par_done_reg367_out;
  wire par_done_reg367_done;
  wire par_done_reg368_in;
  wire par_done_reg368_write_en;
  wire par_done_reg368_clk;
  wire par_done_reg368_out;
  wire par_done_reg368_done;
  wire par_reset17_in;
  wire par_reset17_write_en;
  wire par_reset17_clk;
  wire par_reset17_out;
  wire par_reset17_done;
  wire par_done_reg369_in;
  wire par_done_reg369_write_en;
  wire par_done_reg369_clk;
  wire par_done_reg369_out;
  wire par_done_reg369_done;
  wire par_done_reg370_in;
  wire par_done_reg370_write_en;
  wire par_done_reg370_clk;
  wire par_done_reg370_out;
  wire par_done_reg370_done;
  wire par_done_reg371_in;
  wire par_done_reg371_write_en;
  wire par_done_reg371_clk;
  wire par_done_reg371_out;
  wire par_done_reg371_done;
  wire par_done_reg372_in;
  wire par_done_reg372_write_en;
  wire par_done_reg372_clk;
  wire par_done_reg372_out;
  wire par_done_reg372_done;
  wire par_done_reg373_in;
  wire par_done_reg373_write_en;
  wire par_done_reg373_clk;
  wire par_done_reg373_out;
  wire par_done_reg373_done;
  wire par_done_reg374_in;
  wire par_done_reg374_write_en;
  wire par_done_reg374_clk;
  wire par_done_reg374_out;
  wire par_done_reg374_done;
  wire par_done_reg375_in;
  wire par_done_reg375_write_en;
  wire par_done_reg375_clk;
  wire par_done_reg375_out;
  wire par_done_reg375_done;
  wire par_done_reg376_in;
  wire par_done_reg376_write_en;
  wire par_done_reg376_clk;
  wire par_done_reg376_out;
  wire par_done_reg376_done;
  wire par_done_reg377_in;
  wire par_done_reg377_write_en;
  wire par_done_reg377_clk;
  wire par_done_reg377_out;
  wire par_done_reg377_done;
  wire par_done_reg378_in;
  wire par_done_reg378_write_en;
  wire par_done_reg378_clk;
  wire par_done_reg378_out;
  wire par_done_reg378_done;
  wire par_done_reg379_in;
  wire par_done_reg379_write_en;
  wire par_done_reg379_clk;
  wire par_done_reg379_out;
  wire par_done_reg379_done;
  wire par_done_reg380_in;
  wire par_done_reg380_write_en;
  wire par_done_reg380_clk;
  wire par_done_reg380_out;
  wire par_done_reg380_done;
  wire par_done_reg381_in;
  wire par_done_reg381_write_en;
  wire par_done_reg381_clk;
  wire par_done_reg381_out;
  wire par_done_reg381_done;
  wire par_done_reg382_in;
  wire par_done_reg382_write_en;
  wire par_done_reg382_clk;
  wire par_done_reg382_out;
  wire par_done_reg382_done;
  wire par_done_reg383_in;
  wire par_done_reg383_write_en;
  wire par_done_reg383_clk;
  wire par_done_reg383_out;
  wire par_done_reg383_done;
  wire par_done_reg384_in;
  wire par_done_reg384_write_en;
  wire par_done_reg384_clk;
  wire par_done_reg384_out;
  wire par_done_reg384_done;
  wire par_done_reg385_in;
  wire par_done_reg385_write_en;
  wire par_done_reg385_clk;
  wire par_done_reg385_out;
  wire par_done_reg385_done;
  wire par_done_reg386_in;
  wire par_done_reg386_write_en;
  wire par_done_reg386_clk;
  wire par_done_reg386_out;
  wire par_done_reg386_done;
  wire par_done_reg387_in;
  wire par_done_reg387_write_en;
  wire par_done_reg387_clk;
  wire par_done_reg387_out;
  wire par_done_reg387_done;
  wire par_done_reg388_in;
  wire par_done_reg388_write_en;
  wire par_done_reg388_clk;
  wire par_done_reg388_out;
  wire par_done_reg388_done;
  wire par_done_reg389_in;
  wire par_done_reg389_write_en;
  wire par_done_reg389_clk;
  wire par_done_reg389_out;
  wire par_done_reg389_done;
  wire par_done_reg390_in;
  wire par_done_reg390_write_en;
  wire par_done_reg390_clk;
  wire par_done_reg390_out;
  wire par_done_reg390_done;
  wire par_done_reg391_in;
  wire par_done_reg391_write_en;
  wire par_done_reg391_clk;
  wire par_done_reg391_out;
  wire par_done_reg391_done;
  wire par_done_reg392_in;
  wire par_done_reg392_write_en;
  wire par_done_reg392_clk;
  wire par_done_reg392_out;
  wire par_done_reg392_done;
  wire par_done_reg393_in;
  wire par_done_reg393_write_en;
  wire par_done_reg393_clk;
  wire par_done_reg393_out;
  wire par_done_reg393_done;
  wire par_done_reg394_in;
  wire par_done_reg394_write_en;
  wire par_done_reg394_clk;
  wire par_done_reg394_out;
  wire par_done_reg394_done;
  wire par_done_reg395_in;
  wire par_done_reg395_write_en;
  wire par_done_reg395_clk;
  wire par_done_reg395_out;
  wire par_done_reg395_done;
  wire par_done_reg396_in;
  wire par_done_reg396_write_en;
  wire par_done_reg396_clk;
  wire par_done_reg396_out;
  wire par_done_reg396_done;
  wire par_done_reg397_in;
  wire par_done_reg397_write_en;
  wire par_done_reg397_clk;
  wire par_done_reg397_out;
  wire par_done_reg397_done;
  wire par_done_reg398_in;
  wire par_done_reg398_write_en;
  wire par_done_reg398_clk;
  wire par_done_reg398_out;
  wire par_done_reg398_done;
  wire par_done_reg399_in;
  wire par_done_reg399_write_en;
  wire par_done_reg399_clk;
  wire par_done_reg399_out;
  wire par_done_reg399_done;
  wire par_done_reg400_in;
  wire par_done_reg400_write_en;
  wire par_done_reg400_clk;
  wire par_done_reg400_out;
  wire par_done_reg400_done;
  wire par_done_reg401_in;
  wire par_done_reg401_write_en;
  wire par_done_reg401_clk;
  wire par_done_reg401_out;
  wire par_done_reg401_done;
  wire par_reset18_in;
  wire par_reset18_write_en;
  wire par_reset18_clk;
  wire par_reset18_out;
  wire par_reset18_done;
  wire par_done_reg402_in;
  wire par_done_reg402_write_en;
  wire par_done_reg402_clk;
  wire par_done_reg402_out;
  wire par_done_reg402_done;
  wire par_done_reg403_in;
  wire par_done_reg403_write_en;
  wire par_done_reg403_clk;
  wire par_done_reg403_out;
  wire par_done_reg403_done;
  wire par_done_reg404_in;
  wire par_done_reg404_write_en;
  wire par_done_reg404_clk;
  wire par_done_reg404_out;
  wire par_done_reg404_done;
  wire par_done_reg405_in;
  wire par_done_reg405_write_en;
  wire par_done_reg405_clk;
  wire par_done_reg405_out;
  wire par_done_reg405_done;
  wire par_done_reg406_in;
  wire par_done_reg406_write_en;
  wire par_done_reg406_clk;
  wire par_done_reg406_out;
  wire par_done_reg406_done;
  wire par_done_reg407_in;
  wire par_done_reg407_write_en;
  wire par_done_reg407_clk;
  wire par_done_reg407_out;
  wire par_done_reg407_done;
  wire par_done_reg408_in;
  wire par_done_reg408_write_en;
  wire par_done_reg408_clk;
  wire par_done_reg408_out;
  wire par_done_reg408_done;
  wire par_done_reg409_in;
  wire par_done_reg409_write_en;
  wire par_done_reg409_clk;
  wire par_done_reg409_out;
  wire par_done_reg409_done;
  wire par_done_reg410_in;
  wire par_done_reg410_write_en;
  wire par_done_reg410_clk;
  wire par_done_reg410_out;
  wire par_done_reg410_done;
  wire par_done_reg411_in;
  wire par_done_reg411_write_en;
  wire par_done_reg411_clk;
  wire par_done_reg411_out;
  wire par_done_reg411_done;
  wire par_done_reg412_in;
  wire par_done_reg412_write_en;
  wire par_done_reg412_clk;
  wire par_done_reg412_out;
  wire par_done_reg412_done;
  wire par_done_reg413_in;
  wire par_done_reg413_write_en;
  wire par_done_reg413_clk;
  wire par_done_reg413_out;
  wire par_done_reg413_done;
  wire par_done_reg414_in;
  wire par_done_reg414_write_en;
  wire par_done_reg414_clk;
  wire par_done_reg414_out;
  wire par_done_reg414_done;
  wire par_done_reg415_in;
  wire par_done_reg415_write_en;
  wire par_done_reg415_clk;
  wire par_done_reg415_out;
  wire par_done_reg415_done;
  wire par_done_reg416_in;
  wire par_done_reg416_write_en;
  wire par_done_reg416_clk;
  wire par_done_reg416_out;
  wire par_done_reg416_done;
  wire par_done_reg417_in;
  wire par_done_reg417_write_en;
  wire par_done_reg417_clk;
  wire par_done_reg417_out;
  wire par_done_reg417_done;
  wire par_done_reg418_in;
  wire par_done_reg418_write_en;
  wire par_done_reg418_clk;
  wire par_done_reg418_out;
  wire par_done_reg418_done;
  wire par_done_reg419_in;
  wire par_done_reg419_write_en;
  wire par_done_reg419_clk;
  wire par_done_reg419_out;
  wire par_done_reg419_done;
  wire par_done_reg420_in;
  wire par_done_reg420_write_en;
  wire par_done_reg420_clk;
  wire par_done_reg420_out;
  wire par_done_reg420_done;
  wire par_done_reg421_in;
  wire par_done_reg421_write_en;
  wire par_done_reg421_clk;
  wire par_done_reg421_out;
  wire par_done_reg421_done;
  wire par_done_reg422_in;
  wire par_done_reg422_write_en;
  wire par_done_reg422_clk;
  wire par_done_reg422_out;
  wire par_done_reg422_done;
  wire par_done_reg423_in;
  wire par_done_reg423_write_en;
  wire par_done_reg423_clk;
  wire par_done_reg423_out;
  wire par_done_reg423_done;
  wire par_done_reg424_in;
  wire par_done_reg424_write_en;
  wire par_done_reg424_clk;
  wire par_done_reg424_out;
  wire par_done_reg424_done;
  wire par_done_reg425_in;
  wire par_done_reg425_write_en;
  wire par_done_reg425_clk;
  wire par_done_reg425_out;
  wire par_done_reg425_done;
  wire par_done_reg426_in;
  wire par_done_reg426_write_en;
  wire par_done_reg426_clk;
  wire par_done_reg426_out;
  wire par_done_reg426_done;
  wire par_done_reg427_in;
  wire par_done_reg427_write_en;
  wire par_done_reg427_clk;
  wire par_done_reg427_out;
  wire par_done_reg427_done;
  wire par_done_reg428_in;
  wire par_done_reg428_write_en;
  wire par_done_reg428_clk;
  wire par_done_reg428_out;
  wire par_done_reg428_done;
  wire par_done_reg429_in;
  wire par_done_reg429_write_en;
  wire par_done_reg429_clk;
  wire par_done_reg429_out;
  wire par_done_reg429_done;
  wire par_done_reg430_in;
  wire par_done_reg430_write_en;
  wire par_done_reg430_clk;
  wire par_done_reg430_out;
  wire par_done_reg430_done;
  wire par_done_reg431_in;
  wire par_done_reg431_write_en;
  wire par_done_reg431_clk;
  wire par_done_reg431_out;
  wire par_done_reg431_done;
  wire par_done_reg432_in;
  wire par_done_reg432_write_en;
  wire par_done_reg432_clk;
  wire par_done_reg432_out;
  wire par_done_reg432_done;
  wire par_done_reg433_in;
  wire par_done_reg433_write_en;
  wire par_done_reg433_clk;
  wire par_done_reg433_out;
  wire par_done_reg433_done;
  wire par_done_reg434_in;
  wire par_done_reg434_write_en;
  wire par_done_reg434_clk;
  wire par_done_reg434_out;
  wire par_done_reg434_done;
  wire par_done_reg435_in;
  wire par_done_reg435_write_en;
  wire par_done_reg435_clk;
  wire par_done_reg435_out;
  wire par_done_reg435_done;
  wire par_done_reg436_in;
  wire par_done_reg436_write_en;
  wire par_done_reg436_clk;
  wire par_done_reg436_out;
  wire par_done_reg436_done;
  wire par_done_reg437_in;
  wire par_done_reg437_write_en;
  wire par_done_reg437_clk;
  wire par_done_reg437_out;
  wire par_done_reg437_done;
  wire par_done_reg438_in;
  wire par_done_reg438_write_en;
  wire par_done_reg438_clk;
  wire par_done_reg438_out;
  wire par_done_reg438_done;
  wire par_done_reg439_in;
  wire par_done_reg439_write_en;
  wire par_done_reg439_clk;
  wire par_done_reg439_out;
  wire par_done_reg439_done;
  wire par_done_reg440_in;
  wire par_done_reg440_write_en;
  wire par_done_reg440_clk;
  wire par_done_reg440_out;
  wire par_done_reg440_done;
  wire par_done_reg441_in;
  wire par_done_reg441_write_en;
  wire par_done_reg441_clk;
  wire par_done_reg441_out;
  wire par_done_reg441_done;
  wire par_done_reg442_in;
  wire par_done_reg442_write_en;
  wire par_done_reg442_clk;
  wire par_done_reg442_out;
  wire par_done_reg442_done;
  wire par_done_reg443_in;
  wire par_done_reg443_write_en;
  wire par_done_reg443_clk;
  wire par_done_reg443_out;
  wire par_done_reg443_done;
  wire par_done_reg444_in;
  wire par_done_reg444_write_en;
  wire par_done_reg444_clk;
  wire par_done_reg444_out;
  wire par_done_reg444_done;
  wire par_done_reg445_in;
  wire par_done_reg445_write_en;
  wire par_done_reg445_clk;
  wire par_done_reg445_out;
  wire par_done_reg445_done;
  wire par_done_reg446_in;
  wire par_done_reg446_write_en;
  wire par_done_reg446_clk;
  wire par_done_reg446_out;
  wire par_done_reg446_done;
  wire par_done_reg447_in;
  wire par_done_reg447_write_en;
  wire par_done_reg447_clk;
  wire par_done_reg447_out;
  wire par_done_reg447_done;
  wire par_done_reg448_in;
  wire par_done_reg448_write_en;
  wire par_done_reg448_clk;
  wire par_done_reg448_out;
  wire par_done_reg448_done;
  wire par_done_reg449_in;
  wire par_done_reg449_write_en;
  wire par_done_reg449_clk;
  wire par_done_reg449_out;
  wire par_done_reg449_done;
  wire par_done_reg450_in;
  wire par_done_reg450_write_en;
  wire par_done_reg450_clk;
  wire par_done_reg450_out;
  wire par_done_reg450_done;
  wire par_done_reg451_in;
  wire par_done_reg451_write_en;
  wire par_done_reg451_clk;
  wire par_done_reg451_out;
  wire par_done_reg451_done;
  wire par_done_reg452_in;
  wire par_done_reg452_write_en;
  wire par_done_reg452_clk;
  wire par_done_reg452_out;
  wire par_done_reg452_done;
  wire par_done_reg453_in;
  wire par_done_reg453_write_en;
  wire par_done_reg453_clk;
  wire par_done_reg453_out;
  wire par_done_reg453_done;
  wire par_done_reg454_in;
  wire par_done_reg454_write_en;
  wire par_done_reg454_clk;
  wire par_done_reg454_out;
  wire par_done_reg454_done;
  wire par_done_reg455_in;
  wire par_done_reg455_write_en;
  wire par_done_reg455_clk;
  wire par_done_reg455_out;
  wire par_done_reg455_done;
  wire par_reset19_in;
  wire par_reset19_write_en;
  wire par_reset19_clk;
  wire par_reset19_out;
  wire par_reset19_done;
  wire par_done_reg456_in;
  wire par_done_reg456_write_en;
  wire par_done_reg456_clk;
  wire par_done_reg456_out;
  wire par_done_reg456_done;
  wire par_done_reg457_in;
  wire par_done_reg457_write_en;
  wire par_done_reg457_clk;
  wire par_done_reg457_out;
  wire par_done_reg457_done;
  wire par_done_reg458_in;
  wire par_done_reg458_write_en;
  wire par_done_reg458_clk;
  wire par_done_reg458_out;
  wire par_done_reg458_done;
  wire par_done_reg459_in;
  wire par_done_reg459_write_en;
  wire par_done_reg459_clk;
  wire par_done_reg459_out;
  wire par_done_reg459_done;
  wire par_done_reg460_in;
  wire par_done_reg460_write_en;
  wire par_done_reg460_clk;
  wire par_done_reg460_out;
  wire par_done_reg460_done;
  wire par_done_reg461_in;
  wire par_done_reg461_write_en;
  wire par_done_reg461_clk;
  wire par_done_reg461_out;
  wire par_done_reg461_done;
  wire par_done_reg462_in;
  wire par_done_reg462_write_en;
  wire par_done_reg462_clk;
  wire par_done_reg462_out;
  wire par_done_reg462_done;
  wire par_done_reg463_in;
  wire par_done_reg463_write_en;
  wire par_done_reg463_clk;
  wire par_done_reg463_out;
  wire par_done_reg463_done;
  wire par_done_reg464_in;
  wire par_done_reg464_write_en;
  wire par_done_reg464_clk;
  wire par_done_reg464_out;
  wire par_done_reg464_done;
  wire par_done_reg465_in;
  wire par_done_reg465_write_en;
  wire par_done_reg465_clk;
  wire par_done_reg465_out;
  wire par_done_reg465_done;
  wire par_done_reg466_in;
  wire par_done_reg466_write_en;
  wire par_done_reg466_clk;
  wire par_done_reg466_out;
  wire par_done_reg466_done;
  wire par_done_reg467_in;
  wire par_done_reg467_write_en;
  wire par_done_reg467_clk;
  wire par_done_reg467_out;
  wire par_done_reg467_done;
  wire par_done_reg468_in;
  wire par_done_reg468_write_en;
  wire par_done_reg468_clk;
  wire par_done_reg468_out;
  wire par_done_reg468_done;
  wire par_done_reg469_in;
  wire par_done_reg469_write_en;
  wire par_done_reg469_clk;
  wire par_done_reg469_out;
  wire par_done_reg469_done;
  wire par_done_reg470_in;
  wire par_done_reg470_write_en;
  wire par_done_reg470_clk;
  wire par_done_reg470_out;
  wire par_done_reg470_done;
  wire par_done_reg471_in;
  wire par_done_reg471_write_en;
  wire par_done_reg471_clk;
  wire par_done_reg471_out;
  wire par_done_reg471_done;
  wire par_done_reg472_in;
  wire par_done_reg472_write_en;
  wire par_done_reg472_clk;
  wire par_done_reg472_out;
  wire par_done_reg472_done;
  wire par_done_reg473_in;
  wire par_done_reg473_write_en;
  wire par_done_reg473_clk;
  wire par_done_reg473_out;
  wire par_done_reg473_done;
  wire par_done_reg474_in;
  wire par_done_reg474_write_en;
  wire par_done_reg474_clk;
  wire par_done_reg474_out;
  wire par_done_reg474_done;
  wire par_done_reg475_in;
  wire par_done_reg475_write_en;
  wire par_done_reg475_clk;
  wire par_done_reg475_out;
  wire par_done_reg475_done;
  wire par_done_reg476_in;
  wire par_done_reg476_write_en;
  wire par_done_reg476_clk;
  wire par_done_reg476_out;
  wire par_done_reg476_done;
  wire par_done_reg477_in;
  wire par_done_reg477_write_en;
  wire par_done_reg477_clk;
  wire par_done_reg477_out;
  wire par_done_reg477_done;
  wire par_done_reg478_in;
  wire par_done_reg478_write_en;
  wire par_done_reg478_clk;
  wire par_done_reg478_out;
  wire par_done_reg478_done;
  wire par_done_reg479_in;
  wire par_done_reg479_write_en;
  wire par_done_reg479_clk;
  wire par_done_reg479_out;
  wire par_done_reg479_done;
  wire par_done_reg480_in;
  wire par_done_reg480_write_en;
  wire par_done_reg480_clk;
  wire par_done_reg480_out;
  wire par_done_reg480_done;
  wire par_done_reg481_in;
  wire par_done_reg481_write_en;
  wire par_done_reg481_clk;
  wire par_done_reg481_out;
  wire par_done_reg481_done;
  wire par_done_reg482_in;
  wire par_done_reg482_write_en;
  wire par_done_reg482_clk;
  wire par_done_reg482_out;
  wire par_done_reg482_done;
  wire par_done_reg483_in;
  wire par_done_reg483_write_en;
  wire par_done_reg483_clk;
  wire par_done_reg483_out;
  wire par_done_reg483_done;
  wire par_done_reg484_in;
  wire par_done_reg484_write_en;
  wire par_done_reg484_clk;
  wire par_done_reg484_out;
  wire par_done_reg484_done;
  wire par_done_reg485_in;
  wire par_done_reg485_write_en;
  wire par_done_reg485_clk;
  wire par_done_reg485_out;
  wire par_done_reg485_done;
  wire par_done_reg486_in;
  wire par_done_reg486_write_en;
  wire par_done_reg486_clk;
  wire par_done_reg486_out;
  wire par_done_reg486_done;
  wire par_reset20_in;
  wire par_reset20_write_en;
  wire par_reset20_clk;
  wire par_reset20_out;
  wire par_reset20_done;
  wire par_done_reg487_in;
  wire par_done_reg487_write_en;
  wire par_done_reg487_clk;
  wire par_done_reg487_out;
  wire par_done_reg487_done;
  wire par_done_reg488_in;
  wire par_done_reg488_write_en;
  wire par_done_reg488_clk;
  wire par_done_reg488_out;
  wire par_done_reg488_done;
  wire par_done_reg489_in;
  wire par_done_reg489_write_en;
  wire par_done_reg489_clk;
  wire par_done_reg489_out;
  wire par_done_reg489_done;
  wire par_done_reg490_in;
  wire par_done_reg490_write_en;
  wire par_done_reg490_clk;
  wire par_done_reg490_out;
  wire par_done_reg490_done;
  wire par_done_reg491_in;
  wire par_done_reg491_write_en;
  wire par_done_reg491_clk;
  wire par_done_reg491_out;
  wire par_done_reg491_done;
  wire par_done_reg492_in;
  wire par_done_reg492_write_en;
  wire par_done_reg492_clk;
  wire par_done_reg492_out;
  wire par_done_reg492_done;
  wire par_done_reg493_in;
  wire par_done_reg493_write_en;
  wire par_done_reg493_clk;
  wire par_done_reg493_out;
  wire par_done_reg493_done;
  wire par_done_reg494_in;
  wire par_done_reg494_write_en;
  wire par_done_reg494_clk;
  wire par_done_reg494_out;
  wire par_done_reg494_done;
  wire par_done_reg495_in;
  wire par_done_reg495_write_en;
  wire par_done_reg495_clk;
  wire par_done_reg495_out;
  wire par_done_reg495_done;
  wire par_done_reg496_in;
  wire par_done_reg496_write_en;
  wire par_done_reg496_clk;
  wire par_done_reg496_out;
  wire par_done_reg496_done;
  wire par_done_reg497_in;
  wire par_done_reg497_write_en;
  wire par_done_reg497_clk;
  wire par_done_reg497_out;
  wire par_done_reg497_done;
  wire par_done_reg498_in;
  wire par_done_reg498_write_en;
  wire par_done_reg498_clk;
  wire par_done_reg498_out;
  wire par_done_reg498_done;
  wire par_done_reg499_in;
  wire par_done_reg499_write_en;
  wire par_done_reg499_clk;
  wire par_done_reg499_out;
  wire par_done_reg499_done;
  wire par_done_reg500_in;
  wire par_done_reg500_write_en;
  wire par_done_reg500_clk;
  wire par_done_reg500_out;
  wire par_done_reg500_done;
  wire par_done_reg501_in;
  wire par_done_reg501_write_en;
  wire par_done_reg501_clk;
  wire par_done_reg501_out;
  wire par_done_reg501_done;
  wire par_done_reg502_in;
  wire par_done_reg502_write_en;
  wire par_done_reg502_clk;
  wire par_done_reg502_out;
  wire par_done_reg502_done;
  wire par_done_reg503_in;
  wire par_done_reg503_write_en;
  wire par_done_reg503_clk;
  wire par_done_reg503_out;
  wire par_done_reg503_done;
  wire par_done_reg504_in;
  wire par_done_reg504_write_en;
  wire par_done_reg504_clk;
  wire par_done_reg504_out;
  wire par_done_reg504_done;
  wire par_done_reg505_in;
  wire par_done_reg505_write_en;
  wire par_done_reg505_clk;
  wire par_done_reg505_out;
  wire par_done_reg505_done;
  wire par_done_reg506_in;
  wire par_done_reg506_write_en;
  wire par_done_reg506_clk;
  wire par_done_reg506_out;
  wire par_done_reg506_done;
  wire par_done_reg507_in;
  wire par_done_reg507_write_en;
  wire par_done_reg507_clk;
  wire par_done_reg507_out;
  wire par_done_reg507_done;
  wire par_done_reg508_in;
  wire par_done_reg508_write_en;
  wire par_done_reg508_clk;
  wire par_done_reg508_out;
  wire par_done_reg508_done;
  wire par_done_reg509_in;
  wire par_done_reg509_write_en;
  wire par_done_reg509_clk;
  wire par_done_reg509_out;
  wire par_done_reg509_done;
  wire par_done_reg510_in;
  wire par_done_reg510_write_en;
  wire par_done_reg510_clk;
  wire par_done_reg510_out;
  wire par_done_reg510_done;
  wire par_done_reg511_in;
  wire par_done_reg511_write_en;
  wire par_done_reg511_clk;
  wire par_done_reg511_out;
  wire par_done_reg511_done;
  wire par_done_reg512_in;
  wire par_done_reg512_write_en;
  wire par_done_reg512_clk;
  wire par_done_reg512_out;
  wire par_done_reg512_done;
  wire par_done_reg513_in;
  wire par_done_reg513_write_en;
  wire par_done_reg513_clk;
  wire par_done_reg513_out;
  wire par_done_reg513_done;
  wire par_done_reg514_in;
  wire par_done_reg514_write_en;
  wire par_done_reg514_clk;
  wire par_done_reg514_out;
  wire par_done_reg514_done;
  wire par_done_reg515_in;
  wire par_done_reg515_write_en;
  wire par_done_reg515_clk;
  wire par_done_reg515_out;
  wire par_done_reg515_done;
  wire par_done_reg516_in;
  wire par_done_reg516_write_en;
  wire par_done_reg516_clk;
  wire par_done_reg516_out;
  wire par_done_reg516_done;
  wire par_done_reg517_in;
  wire par_done_reg517_write_en;
  wire par_done_reg517_clk;
  wire par_done_reg517_out;
  wire par_done_reg517_done;
  wire par_done_reg518_in;
  wire par_done_reg518_write_en;
  wire par_done_reg518_clk;
  wire par_done_reg518_out;
  wire par_done_reg518_done;
  wire par_done_reg519_in;
  wire par_done_reg519_write_en;
  wire par_done_reg519_clk;
  wire par_done_reg519_out;
  wire par_done_reg519_done;
  wire par_done_reg520_in;
  wire par_done_reg520_write_en;
  wire par_done_reg520_clk;
  wire par_done_reg520_out;
  wire par_done_reg520_done;
  wire par_done_reg521_in;
  wire par_done_reg521_write_en;
  wire par_done_reg521_clk;
  wire par_done_reg521_out;
  wire par_done_reg521_done;
  wire par_done_reg522_in;
  wire par_done_reg522_write_en;
  wire par_done_reg522_clk;
  wire par_done_reg522_out;
  wire par_done_reg522_done;
  wire par_done_reg523_in;
  wire par_done_reg523_write_en;
  wire par_done_reg523_clk;
  wire par_done_reg523_out;
  wire par_done_reg523_done;
  wire par_done_reg524_in;
  wire par_done_reg524_write_en;
  wire par_done_reg524_clk;
  wire par_done_reg524_out;
  wire par_done_reg524_done;
  wire par_done_reg525_in;
  wire par_done_reg525_write_en;
  wire par_done_reg525_clk;
  wire par_done_reg525_out;
  wire par_done_reg525_done;
  wire par_done_reg526_in;
  wire par_done_reg526_write_en;
  wire par_done_reg526_clk;
  wire par_done_reg526_out;
  wire par_done_reg526_done;
  wire par_done_reg527_in;
  wire par_done_reg527_write_en;
  wire par_done_reg527_clk;
  wire par_done_reg527_out;
  wire par_done_reg527_done;
  wire par_done_reg528_in;
  wire par_done_reg528_write_en;
  wire par_done_reg528_clk;
  wire par_done_reg528_out;
  wire par_done_reg528_done;
  wire par_done_reg529_in;
  wire par_done_reg529_write_en;
  wire par_done_reg529_clk;
  wire par_done_reg529_out;
  wire par_done_reg529_done;
  wire par_done_reg530_in;
  wire par_done_reg530_write_en;
  wire par_done_reg530_clk;
  wire par_done_reg530_out;
  wire par_done_reg530_done;
  wire par_done_reg531_in;
  wire par_done_reg531_write_en;
  wire par_done_reg531_clk;
  wire par_done_reg531_out;
  wire par_done_reg531_done;
  wire par_done_reg532_in;
  wire par_done_reg532_write_en;
  wire par_done_reg532_clk;
  wire par_done_reg532_out;
  wire par_done_reg532_done;
  wire par_done_reg533_in;
  wire par_done_reg533_write_en;
  wire par_done_reg533_clk;
  wire par_done_reg533_out;
  wire par_done_reg533_done;
  wire par_done_reg534_in;
  wire par_done_reg534_write_en;
  wire par_done_reg534_clk;
  wire par_done_reg534_out;
  wire par_done_reg534_done;
  wire par_done_reg535_in;
  wire par_done_reg535_write_en;
  wire par_done_reg535_clk;
  wire par_done_reg535_out;
  wire par_done_reg535_done;
  wire par_done_reg536_in;
  wire par_done_reg536_write_en;
  wire par_done_reg536_clk;
  wire par_done_reg536_out;
  wire par_done_reg536_done;
  wire par_reset21_in;
  wire par_reset21_write_en;
  wire par_reset21_clk;
  wire par_reset21_out;
  wire par_reset21_done;
  wire par_done_reg537_in;
  wire par_done_reg537_write_en;
  wire par_done_reg537_clk;
  wire par_done_reg537_out;
  wire par_done_reg537_done;
  wire par_done_reg538_in;
  wire par_done_reg538_write_en;
  wire par_done_reg538_clk;
  wire par_done_reg538_out;
  wire par_done_reg538_done;
  wire par_done_reg539_in;
  wire par_done_reg539_write_en;
  wire par_done_reg539_clk;
  wire par_done_reg539_out;
  wire par_done_reg539_done;
  wire par_done_reg540_in;
  wire par_done_reg540_write_en;
  wire par_done_reg540_clk;
  wire par_done_reg540_out;
  wire par_done_reg540_done;
  wire par_done_reg541_in;
  wire par_done_reg541_write_en;
  wire par_done_reg541_clk;
  wire par_done_reg541_out;
  wire par_done_reg541_done;
  wire par_done_reg542_in;
  wire par_done_reg542_write_en;
  wire par_done_reg542_clk;
  wire par_done_reg542_out;
  wire par_done_reg542_done;
  wire par_done_reg543_in;
  wire par_done_reg543_write_en;
  wire par_done_reg543_clk;
  wire par_done_reg543_out;
  wire par_done_reg543_done;
  wire par_done_reg544_in;
  wire par_done_reg544_write_en;
  wire par_done_reg544_clk;
  wire par_done_reg544_out;
  wire par_done_reg544_done;
  wire par_done_reg545_in;
  wire par_done_reg545_write_en;
  wire par_done_reg545_clk;
  wire par_done_reg545_out;
  wire par_done_reg545_done;
  wire par_done_reg546_in;
  wire par_done_reg546_write_en;
  wire par_done_reg546_clk;
  wire par_done_reg546_out;
  wire par_done_reg546_done;
  wire par_done_reg547_in;
  wire par_done_reg547_write_en;
  wire par_done_reg547_clk;
  wire par_done_reg547_out;
  wire par_done_reg547_done;
  wire par_done_reg548_in;
  wire par_done_reg548_write_en;
  wire par_done_reg548_clk;
  wire par_done_reg548_out;
  wire par_done_reg548_done;
  wire par_done_reg549_in;
  wire par_done_reg549_write_en;
  wire par_done_reg549_clk;
  wire par_done_reg549_out;
  wire par_done_reg549_done;
  wire par_done_reg550_in;
  wire par_done_reg550_write_en;
  wire par_done_reg550_clk;
  wire par_done_reg550_out;
  wire par_done_reg550_done;
  wire par_done_reg551_in;
  wire par_done_reg551_write_en;
  wire par_done_reg551_clk;
  wire par_done_reg551_out;
  wire par_done_reg551_done;
  wire par_done_reg552_in;
  wire par_done_reg552_write_en;
  wire par_done_reg552_clk;
  wire par_done_reg552_out;
  wire par_done_reg552_done;
  wire par_done_reg553_in;
  wire par_done_reg553_write_en;
  wire par_done_reg553_clk;
  wire par_done_reg553_out;
  wire par_done_reg553_done;
  wire par_done_reg554_in;
  wire par_done_reg554_write_en;
  wire par_done_reg554_clk;
  wire par_done_reg554_out;
  wire par_done_reg554_done;
  wire par_done_reg555_in;
  wire par_done_reg555_write_en;
  wire par_done_reg555_clk;
  wire par_done_reg555_out;
  wire par_done_reg555_done;
  wire par_done_reg556_in;
  wire par_done_reg556_write_en;
  wire par_done_reg556_clk;
  wire par_done_reg556_out;
  wire par_done_reg556_done;
  wire par_done_reg557_in;
  wire par_done_reg557_write_en;
  wire par_done_reg557_clk;
  wire par_done_reg557_out;
  wire par_done_reg557_done;
  wire par_done_reg558_in;
  wire par_done_reg558_write_en;
  wire par_done_reg558_clk;
  wire par_done_reg558_out;
  wire par_done_reg558_done;
  wire par_done_reg559_in;
  wire par_done_reg559_write_en;
  wire par_done_reg559_clk;
  wire par_done_reg559_out;
  wire par_done_reg559_done;
  wire par_done_reg560_in;
  wire par_done_reg560_write_en;
  wire par_done_reg560_clk;
  wire par_done_reg560_out;
  wire par_done_reg560_done;
  wire par_done_reg561_in;
  wire par_done_reg561_write_en;
  wire par_done_reg561_clk;
  wire par_done_reg561_out;
  wire par_done_reg561_done;
  wire par_done_reg562_in;
  wire par_done_reg562_write_en;
  wire par_done_reg562_clk;
  wire par_done_reg562_out;
  wire par_done_reg562_done;
  wire par_done_reg563_in;
  wire par_done_reg563_write_en;
  wire par_done_reg563_clk;
  wire par_done_reg563_out;
  wire par_done_reg563_done;
  wire par_reset22_in;
  wire par_reset22_write_en;
  wire par_reset22_clk;
  wire par_reset22_out;
  wire par_reset22_done;
  wire par_done_reg564_in;
  wire par_done_reg564_write_en;
  wire par_done_reg564_clk;
  wire par_done_reg564_out;
  wire par_done_reg564_done;
  wire par_done_reg565_in;
  wire par_done_reg565_write_en;
  wire par_done_reg565_clk;
  wire par_done_reg565_out;
  wire par_done_reg565_done;
  wire par_done_reg566_in;
  wire par_done_reg566_write_en;
  wire par_done_reg566_clk;
  wire par_done_reg566_out;
  wire par_done_reg566_done;
  wire par_done_reg567_in;
  wire par_done_reg567_write_en;
  wire par_done_reg567_clk;
  wire par_done_reg567_out;
  wire par_done_reg567_done;
  wire par_done_reg568_in;
  wire par_done_reg568_write_en;
  wire par_done_reg568_clk;
  wire par_done_reg568_out;
  wire par_done_reg568_done;
  wire par_done_reg569_in;
  wire par_done_reg569_write_en;
  wire par_done_reg569_clk;
  wire par_done_reg569_out;
  wire par_done_reg569_done;
  wire par_done_reg570_in;
  wire par_done_reg570_write_en;
  wire par_done_reg570_clk;
  wire par_done_reg570_out;
  wire par_done_reg570_done;
  wire par_done_reg571_in;
  wire par_done_reg571_write_en;
  wire par_done_reg571_clk;
  wire par_done_reg571_out;
  wire par_done_reg571_done;
  wire par_done_reg572_in;
  wire par_done_reg572_write_en;
  wire par_done_reg572_clk;
  wire par_done_reg572_out;
  wire par_done_reg572_done;
  wire par_done_reg573_in;
  wire par_done_reg573_write_en;
  wire par_done_reg573_clk;
  wire par_done_reg573_out;
  wire par_done_reg573_done;
  wire par_done_reg574_in;
  wire par_done_reg574_write_en;
  wire par_done_reg574_clk;
  wire par_done_reg574_out;
  wire par_done_reg574_done;
  wire par_done_reg575_in;
  wire par_done_reg575_write_en;
  wire par_done_reg575_clk;
  wire par_done_reg575_out;
  wire par_done_reg575_done;
  wire par_done_reg576_in;
  wire par_done_reg576_write_en;
  wire par_done_reg576_clk;
  wire par_done_reg576_out;
  wire par_done_reg576_done;
  wire par_done_reg577_in;
  wire par_done_reg577_write_en;
  wire par_done_reg577_clk;
  wire par_done_reg577_out;
  wire par_done_reg577_done;
  wire par_done_reg578_in;
  wire par_done_reg578_write_en;
  wire par_done_reg578_clk;
  wire par_done_reg578_out;
  wire par_done_reg578_done;
  wire par_done_reg579_in;
  wire par_done_reg579_write_en;
  wire par_done_reg579_clk;
  wire par_done_reg579_out;
  wire par_done_reg579_done;
  wire par_done_reg580_in;
  wire par_done_reg580_write_en;
  wire par_done_reg580_clk;
  wire par_done_reg580_out;
  wire par_done_reg580_done;
  wire par_done_reg581_in;
  wire par_done_reg581_write_en;
  wire par_done_reg581_clk;
  wire par_done_reg581_out;
  wire par_done_reg581_done;
  wire par_done_reg582_in;
  wire par_done_reg582_write_en;
  wire par_done_reg582_clk;
  wire par_done_reg582_out;
  wire par_done_reg582_done;
  wire par_done_reg583_in;
  wire par_done_reg583_write_en;
  wire par_done_reg583_clk;
  wire par_done_reg583_out;
  wire par_done_reg583_done;
  wire par_done_reg584_in;
  wire par_done_reg584_write_en;
  wire par_done_reg584_clk;
  wire par_done_reg584_out;
  wire par_done_reg584_done;
  wire par_done_reg585_in;
  wire par_done_reg585_write_en;
  wire par_done_reg585_clk;
  wire par_done_reg585_out;
  wire par_done_reg585_done;
  wire par_done_reg586_in;
  wire par_done_reg586_write_en;
  wire par_done_reg586_clk;
  wire par_done_reg586_out;
  wire par_done_reg586_done;
  wire par_done_reg587_in;
  wire par_done_reg587_write_en;
  wire par_done_reg587_clk;
  wire par_done_reg587_out;
  wire par_done_reg587_done;
  wire par_done_reg588_in;
  wire par_done_reg588_write_en;
  wire par_done_reg588_clk;
  wire par_done_reg588_out;
  wire par_done_reg588_done;
  wire par_done_reg589_in;
  wire par_done_reg589_write_en;
  wire par_done_reg589_clk;
  wire par_done_reg589_out;
  wire par_done_reg589_done;
  wire par_done_reg590_in;
  wire par_done_reg590_write_en;
  wire par_done_reg590_clk;
  wire par_done_reg590_out;
  wire par_done_reg590_done;
  wire par_done_reg591_in;
  wire par_done_reg591_write_en;
  wire par_done_reg591_clk;
  wire par_done_reg591_out;
  wire par_done_reg591_done;
  wire par_done_reg592_in;
  wire par_done_reg592_write_en;
  wire par_done_reg592_clk;
  wire par_done_reg592_out;
  wire par_done_reg592_done;
  wire par_done_reg593_in;
  wire par_done_reg593_write_en;
  wire par_done_reg593_clk;
  wire par_done_reg593_out;
  wire par_done_reg593_done;
  wire par_done_reg594_in;
  wire par_done_reg594_write_en;
  wire par_done_reg594_clk;
  wire par_done_reg594_out;
  wire par_done_reg594_done;
  wire par_done_reg595_in;
  wire par_done_reg595_write_en;
  wire par_done_reg595_clk;
  wire par_done_reg595_out;
  wire par_done_reg595_done;
  wire par_done_reg596_in;
  wire par_done_reg596_write_en;
  wire par_done_reg596_clk;
  wire par_done_reg596_out;
  wire par_done_reg596_done;
  wire par_done_reg597_in;
  wire par_done_reg597_write_en;
  wire par_done_reg597_clk;
  wire par_done_reg597_out;
  wire par_done_reg597_done;
  wire par_done_reg598_in;
  wire par_done_reg598_write_en;
  wire par_done_reg598_clk;
  wire par_done_reg598_out;
  wire par_done_reg598_done;
  wire par_done_reg599_in;
  wire par_done_reg599_write_en;
  wire par_done_reg599_clk;
  wire par_done_reg599_out;
  wire par_done_reg599_done;
  wire par_done_reg600_in;
  wire par_done_reg600_write_en;
  wire par_done_reg600_clk;
  wire par_done_reg600_out;
  wire par_done_reg600_done;
  wire par_done_reg601_in;
  wire par_done_reg601_write_en;
  wire par_done_reg601_clk;
  wire par_done_reg601_out;
  wire par_done_reg601_done;
  wire par_done_reg602_in;
  wire par_done_reg602_write_en;
  wire par_done_reg602_clk;
  wire par_done_reg602_out;
  wire par_done_reg602_done;
  wire par_done_reg603_in;
  wire par_done_reg603_write_en;
  wire par_done_reg603_clk;
  wire par_done_reg603_out;
  wire par_done_reg603_done;
  wire par_done_reg604_in;
  wire par_done_reg604_write_en;
  wire par_done_reg604_clk;
  wire par_done_reg604_out;
  wire par_done_reg604_done;
  wire par_done_reg605_in;
  wire par_done_reg605_write_en;
  wire par_done_reg605_clk;
  wire par_done_reg605_out;
  wire par_done_reg605_done;
  wire par_reset23_in;
  wire par_reset23_write_en;
  wire par_reset23_clk;
  wire par_reset23_out;
  wire par_reset23_done;
  wire par_done_reg606_in;
  wire par_done_reg606_write_en;
  wire par_done_reg606_clk;
  wire par_done_reg606_out;
  wire par_done_reg606_done;
  wire par_done_reg607_in;
  wire par_done_reg607_write_en;
  wire par_done_reg607_clk;
  wire par_done_reg607_out;
  wire par_done_reg607_done;
  wire par_done_reg608_in;
  wire par_done_reg608_write_en;
  wire par_done_reg608_clk;
  wire par_done_reg608_out;
  wire par_done_reg608_done;
  wire par_done_reg609_in;
  wire par_done_reg609_write_en;
  wire par_done_reg609_clk;
  wire par_done_reg609_out;
  wire par_done_reg609_done;
  wire par_done_reg610_in;
  wire par_done_reg610_write_en;
  wire par_done_reg610_clk;
  wire par_done_reg610_out;
  wire par_done_reg610_done;
  wire par_done_reg611_in;
  wire par_done_reg611_write_en;
  wire par_done_reg611_clk;
  wire par_done_reg611_out;
  wire par_done_reg611_done;
  wire par_done_reg612_in;
  wire par_done_reg612_write_en;
  wire par_done_reg612_clk;
  wire par_done_reg612_out;
  wire par_done_reg612_done;
  wire par_done_reg613_in;
  wire par_done_reg613_write_en;
  wire par_done_reg613_clk;
  wire par_done_reg613_out;
  wire par_done_reg613_done;
  wire par_done_reg614_in;
  wire par_done_reg614_write_en;
  wire par_done_reg614_clk;
  wire par_done_reg614_out;
  wire par_done_reg614_done;
  wire par_done_reg615_in;
  wire par_done_reg615_write_en;
  wire par_done_reg615_clk;
  wire par_done_reg615_out;
  wire par_done_reg615_done;
  wire par_done_reg616_in;
  wire par_done_reg616_write_en;
  wire par_done_reg616_clk;
  wire par_done_reg616_out;
  wire par_done_reg616_done;
  wire par_done_reg617_in;
  wire par_done_reg617_write_en;
  wire par_done_reg617_clk;
  wire par_done_reg617_out;
  wire par_done_reg617_done;
  wire par_done_reg618_in;
  wire par_done_reg618_write_en;
  wire par_done_reg618_clk;
  wire par_done_reg618_out;
  wire par_done_reg618_done;
  wire par_done_reg619_in;
  wire par_done_reg619_write_en;
  wire par_done_reg619_clk;
  wire par_done_reg619_out;
  wire par_done_reg619_done;
  wire par_done_reg620_in;
  wire par_done_reg620_write_en;
  wire par_done_reg620_clk;
  wire par_done_reg620_out;
  wire par_done_reg620_done;
  wire par_done_reg621_in;
  wire par_done_reg621_write_en;
  wire par_done_reg621_clk;
  wire par_done_reg621_out;
  wire par_done_reg621_done;
  wire par_done_reg622_in;
  wire par_done_reg622_write_en;
  wire par_done_reg622_clk;
  wire par_done_reg622_out;
  wire par_done_reg622_done;
  wire par_done_reg623_in;
  wire par_done_reg623_write_en;
  wire par_done_reg623_clk;
  wire par_done_reg623_out;
  wire par_done_reg623_done;
  wire par_done_reg624_in;
  wire par_done_reg624_write_en;
  wire par_done_reg624_clk;
  wire par_done_reg624_out;
  wire par_done_reg624_done;
  wire par_done_reg625_in;
  wire par_done_reg625_write_en;
  wire par_done_reg625_clk;
  wire par_done_reg625_out;
  wire par_done_reg625_done;
  wire par_done_reg626_in;
  wire par_done_reg626_write_en;
  wire par_done_reg626_clk;
  wire par_done_reg626_out;
  wire par_done_reg626_done;
  wire par_reset24_in;
  wire par_reset24_write_en;
  wire par_reset24_clk;
  wire par_reset24_out;
  wire par_reset24_done;
  wire par_done_reg627_in;
  wire par_done_reg627_write_en;
  wire par_done_reg627_clk;
  wire par_done_reg627_out;
  wire par_done_reg627_done;
  wire par_done_reg628_in;
  wire par_done_reg628_write_en;
  wire par_done_reg628_clk;
  wire par_done_reg628_out;
  wire par_done_reg628_done;
  wire par_done_reg629_in;
  wire par_done_reg629_write_en;
  wire par_done_reg629_clk;
  wire par_done_reg629_out;
  wire par_done_reg629_done;
  wire par_done_reg630_in;
  wire par_done_reg630_write_en;
  wire par_done_reg630_clk;
  wire par_done_reg630_out;
  wire par_done_reg630_done;
  wire par_done_reg631_in;
  wire par_done_reg631_write_en;
  wire par_done_reg631_clk;
  wire par_done_reg631_out;
  wire par_done_reg631_done;
  wire par_done_reg632_in;
  wire par_done_reg632_write_en;
  wire par_done_reg632_clk;
  wire par_done_reg632_out;
  wire par_done_reg632_done;
  wire par_done_reg633_in;
  wire par_done_reg633_write_en;
  wire par_done_reg633_clk;
  wire par_done_reg633_out;
  wire par_done_reg633_done;
  wire par_done_reg634_in;
  wire par_done_reg634_write_en;
  wire par_done_reg634_clk;
  wire par_done_reg634_out;
  wire par_done_reg634_done;
  wire par_done_reg635_in;
  wire par_done_reg635_write_en;
  wire par_done_reg635_clk;
  wire par_done_reg635_out;
  wire par_done_reg635_done;
  wire par_done_reg636_in;
  wire par_done_reg636_write_en;
  wire par_done_reg636_clk;
  wire par_done_reg636_out;
  wire par_done_reg636_done;
  wire par_done_reg637_in;
  wire par_done_reg637_write_en;
  wire par_done_reg637_clk;
  wire par_done_reg637_out;
  wire par_done_reg637_done;
  wire par_done_reg638_in;
  wire par_done_reg638_write_en;
  wire par_done_reg638_clk;
  wire par_done_reg638_out;
  wire par_done_reg638_done;
  wire par_done_reg639_in;
  wire par_done_reg639_write_en;
  wire par_done_reg639_clk;
  wire par_done_reg639_out;
  wire par_done_reg639_done;
  wire par_done_reg640_in;
  wire par_done_reg640_write_en;
  wire par_done_reg640_clk;
  wire par_done_reg640_out;
  wire par_done_reg640_done;
  wire par_done_reg641_in;
  wire par_done_reg641_write_en;
  wire par_done_reg641_clk;
  wire par_done_reg641_out;
  wire par_done_reg641_done;
  wire par_done_reg642_in;
  wire par_done_reg642_write_en;
  wire par_done_reg642_clk;
  wire par_done_reg642_out;
  wire par_done_reg642_done;
  wire par_done_reg643_in;
  wire par_done_reg643_write_en;
  wire par_done_reg643_clk;
  wire par_done_reg643_out;
  wire par_done_reg643_done;
  wire par_done_reg644_in;
  wire par_done_reg644_write_en;
  wire par_done_reg644_clk;
  wire par_done_reg644_out;
  wire par_done_reg644_done;
  wire par_done_reg645_in;
  wire par_done_reg645_write_en;
  wire par_done_reg645_clk;
  wire par_done_reg645_out;
  wire par_done_reg645_done;
  wire par_done_reg646_in;
  wire par_done_reg646_write_en;
  wire par_done_reg646_clk;
  wire par_done_reg646_out;
  wire par_done_reg646_done;
  wire par_done_reg647_in;
  wire par_done_reg647_write_en;
  wire par_done_reg647_clk;
  wire par_done_reg647_out;
  wire par_done_reg647_done;
  wire par_done_reg648_in;
  wire par_done_reg648_write_en;
  wire par_done_reg648_clk;
  wire par_done_reg648_out;
  wire par_done_reg648_done;
  wire par_done_reg649_in;
  wire par_done_reg649_write_en;
  wire par_done_reg649_clk;
  wire par_done_reg649_out;
  wire par_done_reg649_done;
  wire par_done_reg650_in;
  wire par_done_reg650_write_en;
  wire par_done_reg650_clk;
  wire par_done_reg650_out;
  wire par_done_reg650_done;
  wire par_done_reg651_in;
  wire par_done_reg651_write_en;
  wire par_done_reg651_clk;
  wire par_done_reg651_out;
  wire par_done_reg651_done;
  wire par_done_reg652_in;
  wire par_done_reg652_write_en;
  wire par_done_reg652_clk;
  wire par_done_reg652_out;
  wire par_done_reg652_done;
  wire par_done_reg653_in;
  wire par_done_reg653_write_en;
  wire par_done_reg653_clk;
  wire par_done_reg653_out;
  wire par_done_reg653_done;
  wire par_done_reg654_in;
  wire par_done_reg654_write_en;
  wire par_done_reg654_clk;
  wire par_done_reg654_out;
  wire par_done_reg654_done;
  wire par_done_reg655_in;
  wire par_done_reg655_write_en;
  wire par_done_reg655_clk;
  wire par_done_reg655_out;
  wire par_done_reg655_done;
  wire par_done_reg656_in;
  wire par_done_reg656_write_en;
  wire par_done_reg656_clk;
  wire par_done_reg656_out;
  wire par_done_reg656_done;
  wire par_reset25_in;
  wire par_reset25_write_en;
  wire par_reset25_clk;
  wire par_reset25_out;
  wire par_reset25_done;
  wire par_done_reg657_in;
  wire par_done_reg657_write_en;
  wire par_done_reg657_clk;
  wire par_done_reg657_out;
  wire par_done_reg657_done;
  wire par_done_reg658_in;
  wire par_done_reg658_write_en;
  wire par_done_reg658_clk;
  wire par_done_reg658_out;
  wire par_done_reg658_done;
  wire par_done_reg659_in;
  wire par_done_reg659_write_en;
  wire par_done_reg659_clk;
  wire par_done_reg659_out;
  wire par_done_reg659_done;
  wire par_done_reg660_in;
  wire par_done_reg660_write_en;
  wire par_done_reg660_clk;
  wire par_done_reg660_out;
  wire par_done_reg660_done;
  wire par_done_reg661_in;
  wire par_done_reg661_write_en;
  wire par_done_reg661_clk;
  wire par_done_reg661_out;
  wire par_done_reg661_done;
  wire par_done_reg662_in;
  wire par_done_reg662_write_en;
  wire par_done_reg662_clk;
  wire par_done_reg662_out;
  wire par_done_reg662_done;
  wire par_done_reg663_in;
  wire par_done_reg663_write_en;
  wire par_done_reg663_clk;
  wire par_done_reg663_out;
  wire par_done_reg663_done;
  wire par_done_reg664_in;
  wire par_done_reg664_write_en;
  wire par_done_reg664_clk;
  wire par_done_reg664_out;
  wire par_done_reg664_done;
  wire par_done_reg665_in;
  wire par_done_reg665_write_en;
  wire par_done_reg665_clk;
  wire par_done_reg665_out;
  wire par_done_reg665_done;
  wire par_done_reg666_in;
  wire par_done_reg666_write_en;
  wire par_done_reg666_clk;
  wire par_done_reg666_out;
  wire par_done_reg666_done;
  wire par_done_reg667_in;
  wire par_done_reg667_write_en;
  wire par_done_reg667_clk;
  wire par_done_reg667_out;
  wire par_done_reg667_done;
  wire par_done_reg668_in;
  wire par_done_reg668_write_en;
  wire par_done_reg668_clk;
  wire par_done_reg668_out;
  wire par_done_reg668_done;
  wire par_done_reg669_in;
  wire par_done_reg669_write_en;
  wire par_done_reg669_clk;
  wire par_done_reg669_out;
  wire par_done_reg669_done;
  wire par_done_reg670_in;
  wire par_done_reg670_write_en;
  wire par_done_reg670_clk;
  wire par_done_reg670_out;
  wire par_done_reg670_done;
  wire par_done_reg671_in;
  wire par_done_reg671_write_en;
  wire par_done_reg671_clk;
  wire par_done_reg671_out;
  wire par_done_reg671_done;
  wire par_reset26_in;
  wire par_reset26_write_en;
  wire par_reset26_clk;
  wire par_reset26_out;
  wire par_reset26_done;
  wire par_done_reg672_in;
  wire par_done_reg672_write_en;
  wire par_done_reg672_clk;
  wire par_done_reg672_out;
  wire par_done_reg672_done;
  wire par_done_reg673_in;
  wire par_done_reg673_write_en;
  wire par_done_reg673_clk;
  wire par_done_reg673_out;
  wire par_done_reg673_done;
  wire par_done_reg674_in;
  wire par_done_reg674_write_en;
  wire par_done_reg674_clk;
  wire par_done_reg674_out;
  wire par_done_reg674_done;
  wire par_done_reg675_in;
  wire par_done_reg675_write_en;
  wire par_done_reg675_clk;
  wire par_done_reg675_out;
  wire par_done_reg675_done;
  wire par_done_reg676_in;
  wire par_done_reg676_write_en;
  wire par_done_reg676_clk;
  wire par_done_reg676_out;
  wire par_done_reg676_done;
  wire par_done_reg677_in;
  wire par_done_reg677_write_en;
  wire par_done_reg677_clk;
  wire par_done_reg677_out;
  wire par_done_reg677_done;
  wire par_done_reg678_in;
  wire par_done_reg678_write_en;
  wire par_done_reg678_clk;
  wire par_done_reg678_out;
  wire par_done_reg678_done;
  wire par_done_reg679_in;
  wire par_done_reg679_write_en;
  wire par_done_reg679_clk;
  wire par_done_reg679_out;
  wire par_done_reg679_done;
  wire par_done_reg680_in;
  wire par_done_reg680_write_en;
  wire par_done_reg680_clk;
  wire par_done_reg680_out;
  wire par_done_reg680_done;
  wire par_done_reg681_in;
  wire par_done_reg681_write_en;
  wire par_done_reg681_clk;
  wire par_done_reg681_out;
  wire par_done_reg681_done;
  wire par_done_reg682_in;
  wire par_done_reg682_write_en;
  wire par_done_reg682_clk;
  wire par_done_reg682_out;
  wire par_done_reg682_done;
  wire par_done_reg683_in;
  wire par_done_reg683_write_en;
  wire par_done_reg683_clk;
  wire par_done_reg683_out;
  wire par_done_reg683_done;
  wire par_done_reg684_in;
  wire par_done_reg684_write_en;
  wire par_done_reg684_clk;
  wire par_done_reg684_out;
  wire par_done_reg684_done;
  wire par_done_reg685_in;
  wire par_done_reg685_write_en;
  wire par_done_reg685_clk;
  wire par_done_reg685_out;
  wire par_done_reg685_done;
  wire par_done_reg686_in;
  wire par_done_reg686_write_en;
  wire par_done_reg686_clk;
  wire par_done_reg686_out;
  wire par_done_reg686_done;
  wire par_done_reg687_in;
  wire par_done_reg687_write_en;
  wire par_done_reg687_clk;
  wire par_done_reg687_out;
  wire par_done_reg687_done;
  wire par_done_reg688_in;
  wire par_done_reg688_write_en;
  wire par_done_reg688_clk;
  wire par_done_reg688_out;
  wire par_done_reg688_done;
  wire par_done_reg689_in;
  wire par_done_reg689_write_en;
  wire par_done_reg689_clk;
  wire par_done_reg689_out;
  wire par_done_reg689_done;
  wire par_done_reg690_in;
  wire par_done_reg690_write_en;
  wire par_done_reg690_clk;
  wire par_done_reg690_out;
  wire par_done_reg690_done;
  wire par_done_reg691_in;
  wire par_done_reg691_write_en;
  wire par_done_reg691_clk;
  wire par_done_reg691_out;
  wire par_done_reg691_done;
  wire par_reset27_in;
  wire par_reset27_write_en;
  wire par_reset27_clk;
  wire par_reset27_out;
  wire par_reset27_done;
  wire par_done_reg692_in;
  wire par_done_reg692_write_en;
  wire par_done_reg692_clk;
  wire par_done_reg692_out;
  wire par_done_reg692_done;
  wire par_done_reg693_in;
  wire par_done_reg693_write_en;
  wire par_done_reg693_clk;
  wire par_done_reg693_out;
  wire par_done_reg693_done;
  wire par_done_reg694_in;
  wire par_done_reg694_write_en;
  wire par_done_reg694_clk;
  wire par_done_reg694_out;
  wire par_done_reg694_done;
  wire par_done_reg695_in;
  wire par_done_reg695_write_en;
  wire par_done_reg695_clk;
  wire par_done_reg695_out;
  wire par_done_reg695_done;
  wire par_done_reg696_in;
  wire par_done_reg696_write_en;
  wire par_done_reg696_clk;
  wire par_done_reg696_out;
  wire par_done_reg696_done;
  wire par_done_reg697_in;
  wire par_done_reg697_write_en;
  wire par_done_reg697_clk;
  wire par_done_reg697_out;
  wire par_done_reg697_done;
  wire par_done_reg698_in;
  wire par_done_reg698_write_en;
  wire par_done_reg698_clk;
  wire par_done_reg698_out;
  wire par_done_reg698_done;
  wire par_done_reg699_in;
  wire par_done_reg699_write_en;
  wire par_done_reg699_clk;
  wire par_done_reg699_out;
  wire par_done_reg699_done;
  wire par_done_reg700_in;
  wire par_done_reg700_write_en;
  wire par_done_reg700_clk;
  wire par_done_reg700_out;
  wire par_done_reg700_done;
  wire par_done_reg701_in;
  wire par_done_reg701_write_en;
  wire par_done_reg701_clk;
  wire par_done_reg701_out;
  wire par_done_reg701_done;
  wire par_reset28_in;
  wire par_reset28_write_en;
  wire par_reset28_clk;
  wire par_reset28_out;
  wire par_reset28_done;
  wire par_done_reg702_in;
  wire par_done_reg702_write_en;
  wire par_done_reg702_clk;
  wire par_done_reg702_out;
  wire par_done_reg702_done;
  wire par_done_reg703_in;
  wire par_done_reg703_write_en;
  wire par_done_reg703_clk;
  wire par_done_reg703_out;
  wire par_done_reg703_done;
  wire par_done_reg704_in;
  wire par_done_reg704_write_en;
  wire par_done_reg704_clk;
  wire par_done_reg704_out;
  wire par_done_reg704_done;
  wire par_done_reg705_in;
  wire par_done_reg705_write_en;
  wire par_done_reg705_clk;
  wire par_done_reg705_out;
  wire par_done_reg705_done;
  wire par_done_reg706_in;
  wire par_done_reg706_write_en;
  wire par_done_reg706_clk;
  wire par_done_reg706_out;
  wire par_done_reg706_done;
  wire par_done_reg707_in;
  wire par_done_reg707_write_en;
  wire par_done_reg707_clk;
  wire par_done_reg707_out;
  wire par_done_reg707_done;
  wire par_done_reg708_in;
  wire par_done_reg708_write_en;
  wire par_done_reg708_clk;
  wire par_done_reg708_out;
  wire par_done_reg708_done;
  wire par_done_reg709_in;
  wire par_done_reg709_write_en;
  wire par_done_reg709_clk;
  wire par_done_reg709_out;
  wire par_done_reg709_done;
  wire par_done_reg710_in;
  wire par_done_reg710_write_en;
  wire par_done_reg710_clk;
  wire par_done_reg710_out;
  wire par_done_reg710_done;
  wire par_done_reg711_in;
  wire par_done_reg711_write_en;
  wire par_done_reg711_clk;
  wire par_done_reg711_out;
  wire par_done_reg711_done;
  wire par_done_reg712_in;
  wire par_done_reg712_write_en;
  wire par_done_reg712_clk;
  wire par_done_reg712_out;
  wire par_done_reg712_done;
  wire par_done_reg713_in;
  wire par_done_reg713_write_en;
  wire par_done_reg713_clk;
  wire par_done_reg713_out;
  wire par_done_reg713_done;
  wire par_reset29_in;
  wire par_reset29_write_en;
  wire par_reset29_clk;
  wire par_reset29_out;
  wire par_reset29_done;
  wire par_done_reg714_in;
  wire par_done_reg714_write_en;
  wire par_done_reg714_clk;
  wire par_done_reg714_out;
  wire par_done_reg714_done;
  wire par_done_reg715_in;
  wire par_done_reg715_write_en;
  wire par_done_reg715_clk;
  wire par_done_reg715_out;
  wire par_done_reg715_done;
  wire par_done_reg716_in;
  wire par_done_reg716_write_en;
  wire par_done_reg716_clk;
  wire par_done_reg716_out;
  wire par_done_reg716_done;
  wire par_done_reg717_in;
  wire par_done_reg717_write_en;
  wire par_done_reg717_clk;
  wire par_done_reg717_out;
  wire par_done_reg717_done;
  wire par_done_reg718_in;
  wire par_done_reg718_write_en;
  wire par_done_reg718_clk;
  wire par_done_reg718_out;
  wire par_done_reg718_done;
  wire par_done_reg719_in;
  wire par_done_reg719_write_en;
  wire par_done_reg719_clk;
  wire par_done_reg719_out;
  wire par_done_reg719_done;
  wire par_reset30_in;
  wire par_reset30_write_en;
  wire par_reset30_clk;
  wire par_reset30_out;
  wire par_reset30_done;
  wire par_done_reg720_in;
  wire par_done_reg720_write_en;
  wire par_done_reg720_clk;
  wire par_done_reg720_out;
  wire par_done_reg720_done;
  wire par_done_reg721_in;
  wire par_done_reg721_write_en;
  wire par_done_reg721_clk;
  wire par_done_reg721_out;
  wire par_done_reg721_done;
  wire par_done_reg722_in;
  wire par_done_reg722_write_en;
  wire par_done_reg722_clk;
  wire par_done_reg722_out;
  wire par_done_reg722_done;
  wire par_done_reg723_in;
  wire par_done_reg723_write_en;
  wire par_done_reg723_clk;
  wire par_done_reg723_out;
  wire par_done_reg723_done;
  wire par_done_reg724_in;
  wire par_done_reg724_write_en;
  wire par_done_reg724_clk;
  wire par_done_reg724_out;
  wire par_done_reg724_done;
  wire par_done_reg725_in;
  wire par_done_reg725_write_en;
  wire par_done_reg725_clk;
  wire par_done_reg725_out;
  wire par_done_reg725_done;
  wire par_reset31_in;
  wire par_reset31_write_en;
  wire par_reset31_clk;
  wire par_reset31_out;
  wire par_reset31_done;
  wire par_done_reg726_in;
  wire par_done_reg726_write_en;
  wire par_done_reg726_clk;
  wire par_done_reg726_out;
  wire par_done_reg726_done;
  wire par_done_reg727_in;
  wire par_done_reg727_write_en;
  wire par_done_reg727_clk;
  wire par_done_reg727_out;
  wire par_done_reg727_done;
  wire par_done_reg728_in;
  wire par_done_reg728_write_en;
  wire par_done_reg728_clk;
  wire par_done_reg728_out;
  wire par_done_reg728_done;
  wire par_reset32_in;
  wire par_reset32_write_en;
  wire par_reset32_clk;
  wire par_reset32_out;
  wire par_reset32_done;
  wire par_done_reg729_in;
  wire par_done_reg729_write_en;
  wire par_done_reg729_clk;
  wire par_done_reg729_out;
  wire par_done_reg729_done;
  wire par_done_reg730_in;
  wire par_done_reg730_write_en;
  wire par_done_reg730_clk;
  wire par_done_reg730_out;
  wire par_done_reg730_done;
  wire par_reset33_in;
  wire par_reset33_write_en;
  wire par_reset33_clk;
  wire par_reset33_out;
  wire par_reset33_done;
  wire par_done_reg731_in;
  wire par_done_reg731_write_en;
  wire par_done_reg731_clk;
  wire par_done_reg731_out;
  wire par_done_reg731_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_reg #(32) left_55_read (
      .in(left_55_read_in),
      .write_en(left_55_read_write_en),
      .clk(clk),
      .out(left_55_read_out),
      .done(left_55_read_done)
  );
  
  std_reg #(32) top_55_read (
      .in(top_55_read_in),
      .write_en(top_55_read_write_en),
      .clk(clk),
      .out(top_55_read_out),
      .done(top_55_read_done)
  );
  
  mac_pe #() pe_55 (
      .top(pe_55_top),
      .left(pe_55_left),
      .go(pe_55_go),
      .clk(clk),
      .down(pe_55_down),
      .right(pe_55_right),
      .out(pe_55_out),
      .done(pe_55_done)
  );
  
  std_reg #(32) right_54_write (
      .in(right_54_write_in),
      .write_en(right_54_write_write_en),
      .clk(clk),
      .out(right_54_write_out),
      .done(right_54_write_done)
  );
  
  std_reg #(32) left_54_read (
      .in(left_54_read_in),
      .write_en(left_54_read_write_en),
      .clk(clk),
      .out(left_54_read_out),
      .done(left_54_read_done)
  );
  
  std_reg #(32) top_54_read (
      .in(top_54_read_in),
      .write_en(top_54_read_write_en),
      .clk(clk),
      .out(top_54_read_out),
      .done(top_54_read_done)
  );
  
  mac_pe #() pe_54 (
      .top(pe_54_top),
      .left(pe_54_left),
      .go(pe_54_go),
      .clk(clk),
      .down(pe_54_down),
      .right(pe_54_right),
      .out(pe_54_out),
      .done(pe_54_done)
  );
  
  std_reg #(32) right_53_write (
      .in(right_53_write_in),
      .write_en(right_53_write_write_en),
      .clk(clk),
      .out(right_53_write_out),
      .done(right_53_write_done)
  );
  
  std_reg #(32) left_53_read (
      .in(left_53_read_in),
      .write_en(left_53_read_write_en),
      .clk(clk),
      .out(left_53_read_out),
      .done(left_53_read_done)
  );
  
  std_reg #(32) top_53_read (
      .in(top_53_read_in),
      .write_en(top_53_read_write_en),
      .clk(clk),
      .out(top_53_read_out),
      .done(top_53_read_done)
  );
  
  mac_pe #() pe_53 (
      .top(pe_53_top),
      .left(pe_53_left),
      .go(pe_53_go),
      .clk(clk),
      .down(pe_53_down),
      .right(pe_53_right),
      .out(pe_53_out),
      .done(pe_53_done)
  );
  
  std_reg #(32) right_52_write (
      .in(right_52_write_in),
      .write_en(right_52_write_write_en),
      .clk(clk),
      .out(right_52_write_out),
      .done(right_52_write_done)
  );
  
  std_reg #(32) left_52_read (
      .in(left_52_read_in),
      .write_en(left_52_read_write_en),
      .clk(clk),
      .out(left_52_read_out),
      .done(left_52_read_done)
  );
  
  std_reg #(32) top_52_read (
      .in(top_52_read_in),
      .write_en(top_52_read_write_en),
      .clk(clk),
      .out(top_52_read_out),
      .done(top_52_read_done)
  );
  
  mac_pe #() pe_52 (
      .top(pe_52_top),
      .left(pe_52_left),
      .go(pe_52_go),
      .clk(clk),
      .down(pe_52_down),
      .right(pe_52_right),
      .out(pe_52_out),
      .done(pe_52_done)
  );
  
  std_reg #(32) right_51_write (
      .in(right_51_write_in),
      .write_en(right_51_write_write_en),
      .clk(clk),
      .out(right_51_write_out),
      .done(right_51_write_done)
  );
  
  std_reg #(32) left_51_read (
      .in(left_51_read_in),
      .write_en(left_51_read_write_en),
      .clk(clk),
      .out(left_51_read_out),
      .done(left_51_read_done)
  );
  
  std_reg #(32) top_51_read (
      .in(top_51_read_in),
      .write_en(top_51_read_write_en),
      .clk(clk),
      .out(top_51_read_out),
      .done(top_51_read_done)
  );
  
  mac_pe #() pe_51 (
      .top(pe_51_top),
      .left(pe_51_left),
      .go(pe_51_go),
      .clk(clk),
      .down(pe_51_down),
      .right(pe_51_right),
      .out(pe_51_out),
      .done(pe_51_done)
  );
  
  std_reg #(32) right_50_write (
      .in(right_50_write_in),
      .write_en(right_50_write_write_en),
      .clk(clk),
      .out(right_50_write_out),
      .done(right_50_write_done)
  );
  
  std_reg #(32) left_50_read (
      .in(left_50_read_in),
      .write_en(left_50_read_write_en),
      .clk(clk),
      .out(left_50_read_out),
      .done(left_50_read_done)
  );
  
  std_reg #(32) top_50_read (
      .in(top_50_read_in),
      .write_en(top_50_read_write_en),
      .clk(clk),
      .out(top_50_read_out),
      .done(top_50_read_done)
  );
  
  mac_pe #() pe_50 (
      .top(pe_50_top),
      .left(pe_50_left),
      .go(pe_50_go),
      .clk(clk),
      .down(pe_50_down),
      .right(pe_50_right),
      .out(pe_50_out),
      .done(pe_50_done)
  );
  
  std_reg #(32) down_45_write (
      .in(down_45_write_in),
      .write_en(down_45_write_write_en),
      .clk(clk),
      .out(down_45_write_out),
      .done(down_45_write_done)
  );
  
  std_reg #(32) left_45_read (
      .in(left_45_read_in),
      .write_en(left_45_read_write_en),
      .clk(clk),
      .out(left_45_read_out),
      .done(left_45_read_done)
  );
  
  std_reg #(32) top_45_read (
      .in(top_45_read_in),
      .write_en(top_45_read_write_en),
      .clk(clk),
      .out(top_45_read_out),
      .done(top_45_read_done)
  );
  
  mac_pe #() pe_45 (
      .top(pe_45_top),
      .left(pe_45_left),
      .go(pe_45_go),
      .clk(clk),
      .down(pe_45_down),
      .right(pe_45_right),
      .out(pe_45_out),
      .done(pe_45_done)
  );
  
  std_reg #(32) down_44_write (
      .in(down_44_write_in),
      .write_en(down_44_write_write_en),
      .clk(clk),
      .out(down_44_write_out),
      .done(down_44_write_done)
  );
  
  std_reg #(32) right_44_write (
      .in(right_44_write_in),
      .write_en(right_44_write_write_en),
      .clk(clk),
      .out(right_44_write_out),
      .done(right_44_write_done)
  );
  
  std_reg #(32) left_44_read (
      .in(left_44_read_in),
      .write_en(left_44_read_write_en),
      .clk(clk),
      .out(left_44_read_out),
      .done(left_44_read_done)
  );
  
  std_reg #(32) top_44_read (
      .in(top_44_read_in),
      .write_en(top_44_read_write_en),
      .clk(clk),
      .out(top_44_read_out),
      .done(top_44_read_done)
  );
  
  mac_pe #() pe_44 (
      .top(pe_44_top),
      .left(pe_44_left),
      .go(pe_44_go),
      .clk(clk),
      .down(pe_44_down),
      .right(pe_44_right),
      .out(pe_44_out),
      .done(pe_44_done)
  );
  
  std_reg #(32) down_43_write (
      .in(down_43_write_in),
      .write_en(down_43_write_write_en),
      .clk(clk),
      .out(down_43_write_out),
      .done(down_43_write_done)
  );
  
  std_reg #(32) right_43_write (
      .in(right_43_write_in),
      .write_en(right_43_write_write_en),
      .clk(clk),
      .out(right_43_write_out),
      .done(right_43_write_done)
  );
  
  std_reg #(32) left_43_read (
      .in(left_43_read_in),
      .write_en(left_43_read_write_en),
      .clk(clk),
      .out(left_43_read_out),
      .done(left_43_read_done)
  );
  
  std_reg #(32) top_43_read (
      .in(top_43_read_in),
      .write_en(top_43_read_write_en),
      .clk(clk),
      .out(top_43_read_out),
      .done(top_43_read_done)
  );
  
  mac_pe #() pe_43 (
      .top(pe_43_top),
      .left(pe_43_left),
      .go(pe_43_go),
      .clk(clk),
      .down(pe_43_down),
      .right(pe_43_right),
      .out(pe_43_out),
      .done(pe_43_done)
  );
  
  std_reg #(32) down_42_write (
      .in(down_42_write_in),
      .write_en(down_42_write_write_en),
      .clk(clk),
      .out(down_42_write_out),
      .done(down_42_write_done)
  );
  
  std_reg #(32) right_42_write (
      .in(right_42_write_in),
      .write_en(right_42_write_write_en),
      .clk(clk),
      .out(right_42_write_out),
      .done(right_42_write_done)
  );
  
  std_reg #(32) left_42_read (
      .in(left_42_read_in),
      .write_en(left_42_read_write_en),
      .clk(clk),
      .out(left_42_read_out),
      .done(left_42_read_done)
  );
  
  std_reg #(32) top_42_read (
      .in(top_42_read_in),
      .write_en(top_42_read_write_en),
      .clk(clk),
      .out(top_42_read_out),
      .done(top_42_read_done)
  );
  
  mac_pe #() pe_42 (
      .top(pe_42_top),
      .left(pe_42_left),
      .go(pe_42_go),
      .clk(clk),
      .down(pe_42_down),
      .right(pe_42_right),
      .out(pe_42_out),
      .done(pe_42_done)
  );
  
  std_reg #(32) down_41_write (
      .in(down_41_write_in),
      .write_en(down_41_write_write_en),
      .clk(clk),
      .out(down_41_write_out),
      .done(down_41_write_done)
  );
  
  std_reg #(32) right_41_write (
      .in(right_41_write_in),
      .write_en(right_41_write_write_en),
      .clk(clk),
      .out(right_41_write_out),
      .done(right_41_write_done)
  );
  
  std_reg #(32) left_41_read (
      .in(left_41_read_in),
      .write_en(left_41_read_write_en),
      .clk(clk),
      .out(left_41_read_out),
      .done(left_41_read_done)
  );
  
  std_reg #(32) top_41_read (
      .in(top_41_read_in),
      .write_en(top_41_read_write_en),
      .clk(clk),
      .out(top_41_read_out),
      .done(top_41_read_done)
  );
  
  mac_pe #() pe_41 (
      .top(pe_41_top),
      .left(pe_41_left),
      .go(pe_41_go),
      .clk(clk),
      .down(pe_41_down),
      .right(pe_41_right),
      .out(pe_41_out),
      .done(pe_41_done)
  );
  
  std_reg #(32) down_40_write (
      .in(down_40_write_in),
      .write_en(down_40_write_write_en),
      .clk(clk),
      .out(down_40_write_out),
      .done(down_40_write_done)
  );
  
  std_reg #(32) right_40_write (
      .in(right_40_write_in),
      .write_en(right_40_write_write_en),
      .clk(clk),
      .out(right_40_write_out),
      .done(right_40_write_done)
  );
  
  std_reg #(32) left_40_read (
      .in(left_40_read_in),
      .write_en(left_40_read_write_en),
      .clk(clk),
      .out(left_40_read_out),
      .done(left_40_read_done)
  );
  
  std_reg #(32) top_40_read (
      .in(top_40_read_in),
      .write_en(top_40_read_write_en),
      .clk(clk),
      .out(top_40_read_out),
      .done(top_40_read_done)
  );
  
  mac_pe #() pe_40 (
      .top(pe_40_top),
      .left(pe_40_left),
      .go(pe_40_go),
      .clk(clk),
      .down(pe_40_down),
      .right(pe_40_right),
      .out(pe_40_out),
      .done(pe_40_done)
  );
  
  std_reg #(32) down_35_write (
      .in(down_35_write_in),
      .write_en(down_35_write_write_en),
      .clk(clk),
      .out(down_35_write_out),
      .done(down_35_write_done)
  );
  
  std_reg #(32) left_35_read (
      .in(left_35_read_in),
      .write_en(left_35_read_write_en),
      .clk(clk),
      .out(left_35_read_out),
      .done(left_35_read_done)
  );
  
  std_reg #(32) top_35_read (
      .in(top_35_read_in),
      .write_en(top_35_read_write_en),
      .clk(clk),
      .out(top_35_read_out),
      .done(top_35_read_done)
  );
  
  mac_pe #() pe_35 (
      .top(pe_35_top),
      .left(pe_35_left),
      .go(pe_35_go),
      .clk(clk),
      .down(pe_35_down),
      .right(pe_35_right),
      .out(pe_35_out),
      .done(pe_35_done)
  );
  
  std_reg #(32) down_34_write (
      .in(down_34_write_in),
      .write_en(down_34_write_write_en),
      .clk(clk),
      .out(down_34_write_out),
      .done(down_34_write_done)
  );
  
  std_reg #(32) right_34_write (
      .in(right_34_write_in),
      .write_en(right_34_write_write_en),
      .clk(clk),
      .out(right_34_write_out),
      .done(right_34_write_done)
  );
  
  std_reg #(32) left_34_read (
      .in(left_34_read_in),
      .write_en(left_34_read_write_en),
      .clk(clk),
      .out(left_34_read_out),
      .done(left_34_read_done)
  );
  
  std_reg #(32) top_34_read (
      .in(top_34_read_in),
      .write_en(top_34_read_write_en),
      .clk(clk),
      .out(top_34_read_out),
      .done(top_34_read_done)
  );
  
  mac_pe #() pe_34 (
      .top(pe_34_top),
      .left(pe_34_left),
      .go(pe_34_go),
      .clk(clk),
      .down(pe_34_down),
      .right(pe_34_right),
      .out(pe_34_out),
      .done(pe_34_done)
  );
  
  std_reg #(32) down_33_write (
      .in(down_33_write_in),
      .write_en(down_33_write_write_en),
      .clk(clk),
      .out(down_33_write_out),
      .done(down_33_write_done)
  );
  
  std_reg #(32) right_33_write (
      .in(right_33_write_in),
      .write_en(right_33_write_write_en),
      .clk(clk),
      .out(right_33_write_out),
      .done(right_33_write_done)
  );
  
  std_reg #(32) left_33_read (
      .in(left_33_read_in),
      .write_en(left_33_read_write_en),
      .clk(clk),
      .out(left_33_read_out),
      .done(left_33_read_done)
  );
  
  std_reg #(32) top_33_read (
      .in(top_33_read_in),
      .write_en(top_33_read_write_en),
      .clk(clk),
      .out(top_33_read_out),
      .done(top_33_read_done)
  );
  
  mac_pe #() pe_33 (
      .top(pe_33_top),
      .left(pe_33_left),
      .go(pe_33_go),
      .clk(clk),
      .down(pe_33_down),
      .right(pe_33_right),
      .out(pe_33_out),
      .done(pe_33_done)
  );
  
  std_reg #(32) down_32_write (
      .in(down_32_write_in),
      .write_en(down_32_write_write_en),
      .clk(clk),
      .out(down_32_write_out),
      .done(down_32_write_done)
  );
  
  std_reg #(32) right_32_write (
      .in(right_32_write_in),
      .write_en(right_32_write_write_en),
      .clk(clk),
      .out(right_32_write_out),
      .done(right_32_write_done)
  );
  
  std_reg #(32) left_32_read (
      .in(left_32_read_in),
      .write_en(left_32_read_write_en),
      .clk(clk),
      .out(left_32_read_out),
      .done(left_32_read_done)
  );
  
  std_reg #(32) top_32_read (
      .in(top_32_read_in),
      .write_en(top_32_read_write_en),
      .clk(clk),
      .out(top_32_read_out),
      .done(top_32_read_done)
  );
  
  mac_pe #() pe_32 (
      .top(pe_32_top),
      .left(pe_32_left),
      .go(pe_32_go),
      .clk(clk),
      .down(pe_32_down),
      .right(pe_32_right),
      .out(pe_32_out),
      .done(pe_32_done)
  );
  
  std_reg #(32) down_31_write (
      .in(down_31_write_in),
      .write_en(down_31_write_write_en),
      .clk(clk),
      .out(down_31_write_out),
      .done(down_31_write_done)
  );
  
  std_reg #(32) right_31_write (
      .in(right_31_write_in),
      .write_en(right_31_write_write_en),
      .clk(clk),
      .out(right_31_write_out),
      .done(right_31_write_done)
  );
  
  std_reg #(32) left_31_read (
      .in(left_31_read_in),
      .write_en(left_31_read_write_en),
      .clk(clk),
      .out(left_31_read_out),
      .done(left_31_read_done)
  );
  
  std_reg #(32) top_31_read (
      .in(top_31_read_in),
      .write_en(top_31_read_write_en),
      .clk(clk),
      .out(top_31_read_out),
      .done(top_31_read_done)
  );
  
  mac_pe #() pe_31 (
      .top(pe_31_top),
      .left(pe_31_left),
      .go(pe_31_go),
      .clk(clk),
      .down(pe_31_down),
      .right(pe_31_right),
      .out(pe_31_out),
      .done(pe_31_done)
  );
  
  std_reg #(32) down_30_write (
      .in(down_30_write_in),
      .write_en(down_30_write_write_en),
      .clk(clk),
      .out(down_30_write_out),
      .done(down_30_write_done)
  );
  
  std_reg #(32) right_30_write (
      .in(right_30_write_in),
      .write_en(right_30_write_write_en),
      .clk(clk),
      .out(right_30_write_out),
      .done(right_30_write_done)
  );
  
  std_reg #(32) left_30_read (
      .in(left_30_read_in),
      .write_en(left_30_read_write_en),
      .clk(clk),
      .out(left_30_read_out),
      .done(left_30_read_done)
  );
  
  std_reg #(32) top_30_read (
      .in(top_30_read_in),
      .write_en(top_30_read_write_en),
      .clk(clk),
      .out(top_30_read_out),
      .done(top_30_read_done)
  );
  
  mac_pe #() pe_30 (
      .top(pe_30_top),
      .left(pe_30_left),
      .go(pe_30_go),
      .clk(clk),
      .down(pe_30_down),
      .right(pe_30_right),
      .out(pe_30_out),
      .done(pe_30_done)
  );
  
  std_reg #(32) down_25_write (
      .in(down_25_write_in),
      .write_en(down_25_write_write_en),
      .clk(clk),
      .out(down_25_write_out),
      .done(down_25_write_done)
  );
  
  std_reg #(32) left_25_read (
      .in(left_25_read_in),
      .write_en(left_25_read_write_en),
      .clk(clk),
      .out(left_25_read_out),
      .done(left_25_read_done)
  );
  
  std_reg #(32) top_25_read (
      .in(top_25_read_in),
      .write_en(top_25_read_write_en),
      .clk(clk),
      .out(top_25_read_out),
      .done(top_25_read_done)
  );
  
  mac_pe #() pe_25 (
      .top(pe_25_top),
      .left(pe_25_left),
      .go(pe_25_go),
      .clk(clk),
      .down(pe_25_down),
      .right(pe_25_right),
      .out(pe_25_out),
      .done(pe_25_done)
  );
  
  std_reg #(32) down_24_write (
      .in(down_24_write_in),
      .write_en(down_24_write_write_en),
      .clk(clk),
      .out(down_24_write_out),
      .done(down_24_write_done)
  );
  
  std_reg #(32) right_24_write (
      .in(right_24_write_in),
      .write_en(right_24_write_write_en),
      .clk(clk),
      .out(right_24_write_out),
      .done(right_24_write_done)
  );
  
  std_reg #(32) left_24_read (
      .in(left_24_read_in),
      .write_en(left_24_read_write_en),
      .clk(clk),
      .out(left_24_read_out),
      .done(left_24_read_done)
  );
  
  std_reg #(32) top_24_read (
      .in(top_24_read_in),
      .write_en(top_24_read_write_en),
      .clk(clk),
      .out(top_24_read_out),
      .done(top_24_read_done)
  );
  
  mac_pe #() pe_24 (
      .top(pe_24_top),
      .left(pe_24_left),
      .go(pe_24_go),
      .clk(clk),
      .down(pe_24_down),
      .right(pe_24_right),
      .out(pe_24_out),
      .done(pe_24_done)
  );
  
  std_reg #(32) down_23_write (
      .in(down_23_write_in),
      .write_en(down_23_write_write_en),
      .clk(clk),
      .out(down_23_write_out),
      .done(down_23_write_done)
  );
  
  std_reg #(32) right_23_write (
      .in(right_23_write_in),
      .write_en(right_23_write_write_en),
      .clk(clk),
      .out(right_23_write_out),
      .done(right_23_write_done)
  );
  
  std_reg #(32) left_23_read (
      .in(left_23_read_in),
      .write_en(left_23_read_write_en),
      .clk(clk),
      .out(left_23_read_out),
      .done(left_23_read_done)
  );
  
  std_reg #(32) top_23_read (
      .in(top_23_read_in),
      .write_en(top_23_read_write_en),
      .clk(clk),
      .out(top_23_read_out),
      .done(top_23_read_done)
  );
  
  mac_pe #() pe_23 (
      .top(pe_23_top),
      .left(pe_23_left),
      .go(pe_23_go),
      .clk(clk),
      .down(pe_23_down),
      .right(pe_23_right),
      .out(pe_23_out),
      .done(pe_23_done)
  );
  
  std_reg #(32) down_22_write (
      .in(down_22_write_in),
      .write_en(down_22_write_write_en),
      .clk(clk),
      .out(down_22_write_out),
      .done(down_22_write_done)
  );
  
  std_reg #(32) right_22_write (
      .in(right_22_write_in),
      .write_en(right_22_write_write_en),
      .clk(clk),
      .out(right_22_write_out),
      .done(right_22_write_done)
  );
  
  std_reg #(32) left_22_read (
      .in(left_22_read_in),
      .write_en(left_22_read_write_en),
      .clk(clk),
      .out(left_22_read_out),
      .done(left_22_read_done)
  );
  
  std_reg #(32) top_22_read (
      .in(top_22_read_in),
      .write_en(top_22_read_write_en),
      .clk(clk),
      .out(top_22_read_out),
      .done(top_22_read_done)
  );
  
  mac_pe #() pe_22 (
      .top(pe_22_top),
      .left(pe_22_left),
      .go(pe_22_go),
      .clk(clk),
      .down(pe_22_down),
      .right(pe_22_right),
      .out(pe_22_out),
      .done(pe_22_done)
  );
  
  std_reg #(32) down_21_write (
      .in(down_21_write_in),
      .write_en(down_21_write_write_en),
      .clk(clk),
      .out(down_21_write_out),
      .done(down_21_write_done)
  );
  
  std_reg #(32) right_21_write (
      .in(right_21_write_in),
      .write_en(right_21_write_write_en),
      .clk(clk),
      .out(right_21_write_out),
      .done(right_21_write_done)
  );
  
  std_reg #(32) left_21_read (
      .in(left_21_read_in),
      .write_en(left_21_read_write_en),
      .clk(clk),
      .out(left_21_read_out),
      .done(left_21_read_done)
  );
  
  std_reg #(32) top_21_read (
      .in(top_21_read_in),
      .write_en(top_21_read_write_en),
      .clk(clk),
      .out(top_21_read_out),
      .done(top_21_read_done)
  );
  
  mac_pe #() pe_21 (
      .top(pe_21_top),
      .left(pe_21_left),
      .go(pe_21_go),
      .clk(clk),
      .down(pe_21_down),
      .right(pe_21_right),
      .out(pe_21_out),
      .done(pe_21_done)
  );
  
  std_reg #(32) down_20_write (
      .in(down_20_write_in),
      .write_en(down_20_write_write_en),
      .clk(clk),
      .out(down_20_write_out),
      .done(down_20_write_done)
  );
  
  std_reg #(32) right_20_write (
      .in(right_20_write_in),
      .write_en(right_20_write_write_en),
      .clk(clk),
      .out(right_20_write_out),
      .done(right_20_write_done)
  );
  
  std_reg #(32) left_20_read (
      .in(left_20_read_in),
      .write_en(left_20_read_write_en),
      .clk(clk),
      .out(left_20_read_out),
      .done(left_20_read_done)
  );
  
  std_reg #(32) top_20_read (
      .in(top_20_read_in),
      .write_en(top_20_read_write_en),
      .clk(clk),
      .out(top_20_read_out),
      .done(top_20_read_done)
  );
  
  mac_pe #() pe_20 (
      .top(pe_20_top),
      .left(pe_20_left),
      .go(pe_20_go),
      .clk(clk),
      .down(pe_20_down),
      .right(pe_20_right),
      .out(pe_20_out),
      .done(pe_20_done)
  );
  
  std_reg #(32) down_15_write (
      .in(down_15_write_in),
      .write_en(down_15_write_write_en),
      .clk(clk),
      .out(down_15_write_out),
      .done(down_15_write_done)
  );
  
  std_reg #(32) left_15_read (
      .in(left_15_read_in),
      .write_en(left_15_read_write_en),
      .clk(clk),
      .out(left_15_read_out),
      .done(left_15_read_done)
  );
  
  std_reg #(32) top_15_read (
      .in(top_15_read_in),
      .write_en(top_15_read_write_en),
      .clk(clk),
      .out(top_15_read_out),
      .done(top_15_read_done)
  );
  
  mac_pe #() pe_15 (
      .top(pe_15_top),
      .left(pe_15_left),
      .go(pe_15_go),
      .clk(clk),
      .down(pe_15_down),
      .right(pe_15_right),
      .out(pe_15_out),
      .done(pe_15_done)
  );
  
  std_reg #(32) down_14_write (
      .in(down_14_write_in),
      .write_en(down_14_write_write_en),
      .clk(clk),
      .out(down_14_write_out),
      .done(down_14_write_done)
  );
  
  std_reg #(32) right_14_write (
      .in(right_14_write_in),
      .write_en(right_14_write_write_en),
      .clk(clk),
      .out(right_14_write_out),
      .done(right_14_write_done)
  );
  
  std_reg #(32) left_14_read (
      .in(left_14_read_in),
      .write_en(left_14_read_write_en),
      .clk(clk),
      .out(left_14_read_out),
      .done(left_14_read_done)
  );
  
  std_reg #(32) top_14_read (
      .in(top_14_read_in),
      .write_en(top_14_read_write_en),
      .clk(clk),
      .out(top_14_read_out),
      .done(top_14_read_done)
  );
  
  mac_pe #() pe_14 (
      .top(pe_14_top),
      .left(pe_14_left),
      .go(pe_14_go),
      .clk(clk),
      .down(pe_14_down),
      .right(pe_14_right),
      .out(pe_14_out),
      .done(pe_14_done)
  );
  
  std_reg #(32) down_13_write (
      .in(down_13_write_in),
      .write_en(down_13_write_write_en),
      .clk(clk),
      .out(down_13_write_out),
      .done(down_13_write_done)
  );
  
  std_reg #(32) right_13_write (
      .in(right_13_write_in),
      .write_en(right_13_write_write_en),
      .clk(clk),
      .out(right_13_write_out),
      .done(right_13_write_done)
  );
  
  std_reg #(32) left_13_read (
      .in(left_13_read_in),
      .write_en(left_13_read_write_en),
      .clk(clk),
      .out(left_13_read_out),
      .done(left_13_read_done)
  );
  
  std_reg #(32) top_13_read (
      .in(top_13_read_in),
      .write_en(top_13_read_write_en),
      .clk(clk),
      .out(top_13_read_out),
      .done(top_13_read_done)
  );
  
  mac_pe #() pe_13 (
      .top(pe_13_top),
      .left(pe_13_left),
      .go(pe_13_go),
      .clk(clk),
      .down(pe_13_down),
      .right(pe_13_right),
      .out(pe_13_out),
      .done(pe_13_done)
  );
  
  std_reg #(32) down_12_write (
      .in(down_12_write_in),
      .write_en(down_12_write_write_en),
      .clk(clk),
      .out(down_12_write_out),
      .done(down_12_write_done)
  );
  
  std_reg #(32) right_12_write (
      .in(right_12_write_in),
      .write_en(right_12_write_write_en),
      .clk(clk),
      .out(right_12_write_out),
      .done(right_12_write_done)
  );
  
  std_reg #(32) left_12_read (
      .in(left_12_read_in),
      .write_en(left_12_read_write_en),
      .clk(clk),
      .out(left_12_read_out),
      .done(left_12_read_done)
  );
  
  std_reg #(32) top_12_read (
      .in(top_12_read_in),
      .write_en(top_12_read_write_en),
      .clk(clk),
      .out(top_12_read_out),
      .done(top_12_read_done)
  );
  
  mac_pe #() pe_12 (
      .top(pe_12_top),
      .left(pe_12_left),
      .go(pe_12_go),
      .clk(clk),
      .down(pe_12_down),
      .right(pe_12_right),
      .out(pe_12_out),
      .done(pe_12_done)
  );
  
  std_reg #(32) down_11_write (
      .in(down_11_write_in),
      .write_en(down_11_write_write_en),
      .clk(clk),
      .out(down_11_write_out),
      .done(down_11_write_done)
  );
  
  std_reg #(32) right_11_write (
      .in(right_11_write_in),
      .write_en(right_11_write_write_en),
      .clk(clk),
      .out(right_11_write_out),
      .done(right_11_write_done)
  );
  
  std_reg #(32) left_11_read (
      .in(left_11_read_in),
      .write_en(left_11_read_write_en),
      .clk(clk),
      .out(left_11_read_out),
      .done(left_11_read_done)
  );
  
  std_reg #(32) top_11_read (
      .in(top_11_read_in),
      .write_en(top_11_read_write_en),
      .clk(clk),
      .out(top_11_read_out),
      .done(top_11_read_done)
  );
  
  mac_pe #() pe_11 (
      .top(pe_11_top),
      .left(pe_11_left),
      .go(pe_11_go),
      .clk(clk),
      .down(pe_11_down),
      .right(pe_11_right),
      .out(pe_11_out),
      .done(pe_11_done)
  );
  
  std_reg #(32) down_10_write (
      .in(down_10_write_in),
      .write_en(down_10_write_write_en),
      .clk(clk),
      .out(down_10_write_out),
      .done(down_10_write_done)
  );
  
  std_reg #(32) right_10_write (
      .in(right_10_write_in),
      .write_en(right_10_write_write_en),
      .clk(clk),
      .out(right_10_write_out),
      .done(right_10_write_done)
  );
  
  std_reg #(32) left_10_read (
      .in(left_10_read_in),
      .write_en(left_10_read_write_en),
      .clk(clk),
      .out(left_10_read_out),
      .done(left_10_read_done)
  );
  
  std_reg #(32) top_10_read (
      .in(top_10_read_in),
      .write_en(top_10_read_write_en),
      .clk(clk),
      .out(top_10_read_out),
      .done(top_10_read_done)
  );
  
  mac_pe #() pe_10 (
      .top(pe_10_top),
      .left(pe_10_left),
      .go(pe_10_go),
      .clk(clk),
      .down(pe_10_down),
      .right(pe_10_right),
      .out(pe_10_out),
      .done(pe_10_done)
  );
  
  std_reg #(32) down_05_write (
      .in(down_05_write_in),
      .write_en(down_05_write_write_en),
      .clk(clk),
      .out(down_05_write_out),
      .done(down_05_write_done)
  );
  
  std_reg #(32) left_05_read (
      .in(left_05_read_in),
      .write_en(left_05_read_write_en),
      .clk(clk),
      .out(left_05_read_out),
      .done(left_05_read_done)
  );
  
  std_reg #(32) top_05_read (
      .in(top_05_read_in),
      .write_en(top_05_read_write_en),
      .clk(clk),
      .out(top_05_read_out),
      .done(top_05_read_done)
  );
  
  mac_pe #() pe_05 (
      .top(pe_05_top),
      .left(pe_05_left),
      .go(pe_05_go),
      .clk(clk),
      .down(pe_05_down),
      .right(pe_05_right),
      .out(pe_05_out),
      .done(pe_05_done)
  );
  
  std_reg #(32) down_04_write (
      .in(down_04_write_in),
      .write_en(down_04_write_write_en),
      .clk(clk),
      .out(down_04_write_out),
      .done(down_04_write_done)
  );
  
  std_reg #(32) right_04_write (
      .in(right_04_write_in),
      .write_en(right_04_write_write_en),
      .clk(clk),
      .out(right_04_write_out),
      .done(right_04_write_done)
  );
  
  std_reg #(32) left_04_read (
      .in(left_04_read_in),
      .write_en(left_04_read_write_en),
      .clk(clk),
      .out(left_04_read_out),
      .done(left_04_read_done)
  );
  
  std_reg #(32) top_04_read (
      .in(top_04_read_in),
      .write_en(top_04_read_write_en),
      .clk(clk),
      .out(top_04_read_out),
      .done(top_04_read_done)
  );
  
  mac_pe #() pe_04 (
      .top(pe_04_top),
      .left(pe_04_left),
      .go(pe_04_go),
      .clk(clk),
      .down(pe_04_down),
      .right(pe_04_right),
      .out(pe_04_out),
      .done(pe_04_done)
  );
  
  std_reg #(32) down_03_write (
      .in(down_03_write_in),
      .write_en(down_03_write_write_en),
      .clk(clk),
      .out(down_03_write_out),
      .done(down_03_write_done)
  );
  
  std_reg #(32) right_03_write (
      .in(right_03_write_in),
      .write_en(right_03_write_write_en),
      .clk(clk),
      .out(right_03_write_out),
      .done(right_03_write_done)
  );
  
  std_reg #(32) left_03_read (
      .in(left_03_read_in),
      .write_en(left_03_read_write_en),
      .clk(clk),
      .out(left_03_read_out),
      .done(left_03_read_done)
  );
  
  std_reg #(32) top_03_read (
      .in(top_03_read_in),
      .write_en(top_03_read_write_en),
      .clk(clk),
      .out(top_03_read_out),
      .done(top_03_read_done)
  );
  
  mac_pe #() pe_03 (
      .top(pe_03_top),
      .left(pe_03_left),
      .go(pe_03_go),
      .clk(clk),
      .down(pe_03_down),
      .right(pe_03_right),
      .out(pe_03_out),
      .done(pe_03_done)
  );
  
  std_reg #(32) down_02_write (
      .in(down_02_write_in),
      .write_en(down_02_write_write_en),
      .clk(clk),
      .out(down_02_write_out),
      .done(down_02_write_done)
  );
  
  std_reg #(32) right_02_write (
      .in(right_02_write_in),
      .write_en(right_02_write_write_en),
      .clk(clk),
      .out(right_02_write_out),
      .done(right_02_write_done)
  );
  
  std_reg #(32) left_02_read (
      .in(left_02_read_in),
      .write_en(left_02_read_write_en),
      .clk(clk),
      .out(left_02_read_out),
      .done(left_02_read_done)
  );
  
  std_reg #(32) top_02_read (
      .in(top_02_read_in),
      .write_en(top_02_read_write_en),
      .clk(clk),
      .out(top_02_read_out),
      .done(top_02_read_done)
  );
  
  mac_pe #() pe_02 (
      .top(pe_02_top),
      .left(pe_02_left),
      .go(pe_02_go),
      .clk(clk),
      .down(pe_02_down),
      .right(pe_02_right),
      .out(pe_02_out),
      .done(pe_02_done)
  );
  
  std_reg #(32) down_01_write (
      .in(down_01_write_in),
      .write_en(down_01_write_write_en),
      .clk(clk),
      .out(down_01_write_out),
      .done(down_01_write_done)
  );
  
  std_reg #(32) right_01_write (
      .in(right_01_write_in),
      .write_en(right_01_write_write_en),
      .clk(clk),
      .out(right_01_write_out),
      .done(right_01_write_done)
  );
  
  std_reg #(32) left_01_read (
      .in(left_01_read_in),
      .write_en(left_01_read_write_en),
      .clk(clk),
      .out(left_01_read_out),
      .done(left_01_read_done)
  );
  
  std_reg #(32) top_01_read (
      .in(top_01_read_in),
      .write_en(top_01_read_write_en),
      .clk(clk),
      .out(top_01_read_out),
      .done(top_01_read_done)
  );
  
  mac_pe #() pe_01 (
      .top(pe_01_top),
      .left(pe_01_left),
      .go(pe_01_go),
      .clk(clk),
      .down(pe_01_down),
      .right(pe_01_right),
      .out(pe_01_out),
      .done(pe_01_done)
  );
  
  std_reg #(32) down_00_write (
      .in(down_00_write_in),
      .write_en(down_00_write_write_en),
      .clk(clk),
      .out(down_00_write_out),
      .done(down_00_write_done)
  );
  
  std_reg #(32) right_00_write (
      .in(right_00_write_in),
      .write_en(right_00_write_write_en),
      .clk(clk),
      .out(right_00_write_out),
      .done(right_00_write_done)
  );
  
  std_reg #(32) left_00_read (
      .in(left_00_read_in),
      .write_en(left_00_read_write_en),
      .clk(clk),
      .out(left_00_read_out),
      .done(left_00_read_done)
  );
  
  std_reg #(32) top_00_read (
      .in(top_00_read_in),
      .write_en(top_00_read_write_en),
      .clk(clk),
      .out(top_00_read_out),
      .done(top_00_read_done)
  );
  
  mac_pe #() pe_00 (
      .top(pe_00_top),
      .left(pe_00_left),
      .go(pe_00_go),
      .clk(clk),
      .down(pe_00_down),
      .right(pe_00_right),
      .out(pe_00_out),
      .done(pe_00_done)
  );
  
  std_mem_d1 #(32, 6, 3) l5 (
      .addr0(l5_addr0),
      .write_data(l5_write_data),
      .write_en(l5_write_en),
      .clk(clk),
      .read_data(l5_read_data),
      .done(l5_done)
  );
  
  std_add #(3) l5_add (
      .left(l5_add_left),
      .right(l5_add_right),
      .out(l5_add_out)
  );
  
  std_reg #(3) l5_idx (
      .in(l5_idx_in),
      .write_en(l5_idx_write_en),
      .clk(clk),
      .out(l5_idx_out),
      .done(l5_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) l4 (
      .addr0(l4_addr0),
      .write_data(l4_write_data),
      .write_en(l4_write_en),
      .clk(clk),
      .read_data(l4_read_data),
      .done(l4_done)
  );
  
  std_add #(3) l4_add (
      .left(l4_add_left),
      .right(l4_add_right),
      .out(l4_add_out)
  );
  
  std_reg #(3) l4_idx (
      .in(l4_idx_in),
      .write_en(l4_idx_write_en),
      .clk(clk),
      .out(l4_idx_out),
      .done(l4_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) l3 (
      .addr0(l3_addr0),
      .write_data(l3_write_data),
      .write_en(l3_write_en),
      .clk(clk),
      .read_data(l3_read_data),
      .done(l3_done)
  );
  
  std_add #(3) l3_add (
      .left(l3_add_left),
      .right(l3_add_right),
      .out(l3_add_out)
  );
  
  std_reg #(3) l3_idx (
      .in(l3_idx_in),
      .write_en(l3_idx_write_en),
      .clk(clk),
      .out(l3_idx_out),
      .done(l3_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) l2 (
      .addr0(l2_addr0),
      .write_data(l2_write_data),
      .write_en(l2_write_en),
      .clk(clk),
      .read_data(l2_read_data),
      .done(l2_done)
  );
  
  std_add #(3) l2_add (
      .left(l2_add_left),
      .right(l2_add_right),
      .out(l2_add_out)
  );
  
  std_reg #(3) l2_idx (
      .in(l2_idx_in),
      .write_en(l2_idx_write_en),
      .clk(clk),
      .out(l2_idx_out),
      .done(l2_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) l1 (
      .addr0(l1_addr0),
      .write_data(l1_write_data),
      .write_en(l1_write_en),
      .clk(clk),
      .read_data(l1_read_data),
      .done(l1_done)
  );
  
  std_add #(3) l1_add (
      .left(l1_add_left),
      .right(l1_add_right),
      .out(l1_add_out)
  );
  
  std_reg #(3) l1_idx (
      .in(l1_idx_in),
      .write_en(l1_idx_write_en),
      .clk(clk),
      .out(l1_idx_out),
      .done(l1_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) l0 (
      .addr0(l0_addr0),
      .write_data(l0_write_data),
      .write_en(l0_write_en),
      .clk(clk),
      .read_data(l0_read_data),
      .done(l0_done)
  );
  
  std_add #(3) l0_add (
      .left(l0_add_left),
      .right(l0_add_right),
      .out(l0_add_out)
  );
  
  std_reg #(3) l0_idx (
      .in(l0_idx_in),
      .write_en(l0_idx_write_en),
      .clk(clk),
      .out(l0_idx_out),
      .done(l0_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) t5 (
      .addr0(t5_addr0),
      .write_data(t5_write_data),
      .write_en(t5_write_en),
      .clk(clk),
      .read_data(t5_read_data),
      .done(t5_done)
  );
  
  std_add #(3) t5_add (
      .left(t5_add_left),
      .right(t5_add_right),
      .out(t5_add_out)
  );
  
  std_reg #(3) t5_idx (
      .in(t5_idx_in),
      .write_en(t5_idx_write_en),
      .clk(clk),
      .out(t5_idx_out),
      .done(t5_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) t4 (
      .addr0(t4_addr0),
      .write_data(t4_write_data),
      .write_en(t4_write_en),
      .clk(clk),
      .read_data(t4_read_data),
      .done(t4_done)
  );
  
  std_add #(3) t4_add (
      .left(t4_add_left),
      .right(t4_add_right),
      .out(t4_add_out)
  );
  
  std_reg #(3) t4_idx (
      .in(t4_idx_in),
      .write_en(t4_idx_write_en),
      .clk(clk),
      .out(t4_idx_out),
      .done(t4_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) t3 (
      .addr0(t3_addr0),
      .write_data(t3_write_data),
      .write_en(t3_write_en),
      .clk(clk),
      .read_data(t3_read_data),
      .done(t3_done)
  );
  
  std_add #(3) t3_add (
      .left(t3_add_left),
      .right(t3_add_right),
      .out(t3_add_out)
  );
  
  std_reg #(3) t3_idx (
      .in(t3_idx_in),
      .write_en(t3_idx_write_en),
      .clk(clk),
      .out(t3_idx_out),
      .done(t3_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) t2 (
      .addr0(t2_addr0),
      .write_data(t2_write_data),
      .write_en(t2_write_en),
      .clk(clk),
      .read_data(t2_read_data),
      .done(t2_done)
  );
  
  std_add #(3) t2_add (
      .left(t2_add_left),
      .right(t2_add_right),
      .out(t2_add_out)
  );
  
  std_reg #(3) t2_idx (
      .in(t2_idx_in),
      .write_en(t2_idx_write_en),
      .clk(clk),
      .out(t2_idx_out),
      .done(t2_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) t1 (
      .addr0(t1_addr0),
      .write_data(t1_write_data),
      .write_en(t1_write_en),
      .clk(clk),
      .read_data(t1_read_data),
      .done(t1_done)
  );
  
  std_add #(3) t1_add (
      .left(t1_add_left),
      .right(t1_add_right),
      .out(t1_add_out)
  );
  
  std_reg #(3) t1_idx (
      .in(t1_idx_in),
      .write_en(t1_idx_write_en),
      .clk(clk),
      .out(t1_idx_out),
      .done(t1_idx_done)
  );
  
  std_mem_d1 #(32, 6, 3) t0 (
      .addr0(t0_addr0),
      .write_data(t0_write_data),
      .write_en(t0_write_en),
      .clk(clk),
      .read_data(t0_read_data),
      .done(t0_done)
  );
  
  std_add #(3) t0_add (
      .left(t0_add_left),
      .right(t0_add_right),
      .out(t0_add_out)
  );
  
  std_reg #(3) t0_idx (
      .in(t0_idx_in),
      .write_en(t0_idx_write_en),
      .clk(clk),
      .out(t0_idx_out),
      .done(t0_idx_done)
  );
  
  std_reg #(1) par_reset0 (
      .in(par_reset0_in),
      .write_en(par_reset0_write_en),
      .clk(clk),
      .out(par_reset0_out),
      .done(par_reset0_done)
  );
  
  std_reg #(1) par_done_reg0 (
      .in(par_done_reg0_in),
      .write_en(par_done_reg0_write_en),
      .clk(clk),
      .out(par_done_reg0_out),
      .done(par_done_reg0_done)
  );
  
  std_reg #(1) par_done_reg1 (
      .in(par_done_reg1_in),
      .write_en(par_done_reg1_write_en),
      .clk(clk),
      .out(par_done_reg1_out),
      .done(par_done_reg1_done)
  );
  
  std_reg #(1) par_done_reg2 (
      .in(par_done_reg2_in),
      .write_en(par_done_reg2_write_en),
      .clk(clk),
      .out(par_done_reg2_out),
      .done(par_done_reg2_done)
  );
  
  std_reg #(1) par_done_reg3 (
      .in(par_done_reg3_in),
      .write_en(par_done_reg3_write_en),
      .clk(clk),
      .out(par_done_reg3_out),
      .done(par_done_reg3_done)
  );
  
  std_reg #(1) par_done_reg4 (
      .in(par_done_reg4_in),
      .write_en(par_done_reg4_write_en),
      .clk(clk),
      .out(par_done_reg4_out),
      .done(par_done_reg4_done)
  );
  
  std_reg #(1) par_done_reg5 (
      .in(par_done_reg5_in),
      .write_en(par_done_reg5_write_en),
      .clk(clk),
      .out(par_done_reg5_out),
      .done(par_done_reg5_done)
  );
  
  std_reg #(1) par_done_reg6 (
      .in(par_done_reg6_in),
      .write_en(par_done_reg6_write_en),
      .clk(clk),
      .out(par_done_reg6_out),
      .done(par_done_reg6_done)
  );
  
  std_reg #(1) par_done_reg7 (
      .in(par_done_reg7_in),
      .write_en(par_done_reg7_write_en),
      .clk(clk),
      .out(par_done_reg7_out),
      .done(par_done_reg7_done)
  );
  
  std_reg #(1) par_done_reg8 (
      .in(par_done_reg8_in),
      .write_en(par_done_reg8_write_en),
      .clk(clk),
      .out(par_done_reg8_out),
      .done(par_done_reg8_done)
  );
  
  std_reg #(1) par_done_reg9 (
      .in(par_done_reg9_in),
      .write_en(par_done_reg9_write_en),
      .clk(clk),
      .out(par_done_reg9_out),
      .done(par_done_reg9_done)
  );
  
  std_reg #(1) par_done_reg10 (
      .in(par_done_reg10_in),
      .write_en(par_done_reg10_write_en),
      .clk(clk),
      .out(par_done_reg10_out),
      .done(par_done_reg10_done)
  );
  
  std_reg #(1) par_done_reg11 (
      .in(par_done_reg11_in),
      .write_en(par_done_reg11_write_en),
      .clk(clk),
      .out(par_done_reg11_out),
      .done(par_done_reg11_done)
  );
  
  std_reg #(1) par_reset1 (
      .in(par_reset1_in),
      .write_en(par_reset1_write_en),
      .clk(clk),
      .out(par_reset1_out),
      .done(par_reset1_done)
  );
  
  std_reg #(1) par_done_reg12 (
      .in(par_done_reg12_in),
      .write_en(par_done_reg12_write_en),
      .clk(clk),
      .out(par_done_reg12_out),
      .done(par_done_reg12_done)
  );
  
  std_reg #(1) par_done_reg13 (
      .in(par_done_reg13_in),
      .write_en(par_done_reg13_write_en),
      .clk(clk),
      .out(par_done_reg13_out),
      .done(par_done_reg13_done)
  );
  
  std_reg #(1) par_reset2 (
      .in(par_reset2_in),
      .write_en(par_reset2_write_en),
      .clk(clk),
      .out(par_reset2_out),
      .done(par_reset2_done)
  );
  
  std_reg #(1) par_done_reg14 (
      .in(par_done_reg14_in),
      .write_en(par_done_reg14_write_en),
      .clk(clk),
      .out(par_done_reg14_out),
      .done(par_done_reg14_done)
  );
  
  std_reg #(1) par_done_reg15 (
      .in(par_done_reg15_in),
      .write_en(par_done_reg15_write_en),
      .clk(clk),
      .out(par_done_reg15_out),
      .done(par_done_reg15_done)
  );
  
  std_reg #(1) par_reset3 (
      .in(par_reset3_in),
      .write_en(par_reset3_write_en),
      .clk(clk),
      .out(par_reset3_out),
      .done(par_reset3_done)
  );
  
  std_reg #(1) par_done_reg16 (
      .in(par_done_reg16_in),
      .write_en(par_done_reg16_write_en),
      .clk(clk),
      .out(par_done_reg16_out),
      .done(par_done_reg16_done)
  );
  
  std_reg #(1) par_done_reg17 (
      .in(par_done_reg17_in),
      .write_en(par_done_reg17_write_en),
      .clk(clk),
      .out(par_done_reg17_out),
      .done(par_done_reg17_done)
  );
  
  std_reg #(1) par_done_reg18 (
      .in(par_done_reg18_in),
      .write_en(par_done_reg18_write_en),
      .clk(clk),
      .out(par_done_reg18_out),
      .done(par_done_reg18_done)
  );
  
  std_reg #(1) par_done_reg19 (
      .in(par_done_reg19_in),
      .write_en(par_done_reg19_write_en),
      .clk(clk),
      .out(par_done_reg19_out),
      .done(par_done_reg19_done)
  );
  
  std_reg #(1) par_done_reg20 (
      .in(par_done_reg20_in),
      .write_en(par_done_reg20_write_en),
      .clk(clk),
      .out(par_done_reg20_out),
      .done(par_done_reg20_done)
  );
  
  std_reg #(1) par_reset4 (
      .in(par_reset4_in),
      .write_en(par_reset4_write_en),
      .clk(clk),
      .out(par_reset4_out),
      .done(par_reset4_done)
  );
  
  std_reg #(1) par_done_reg21 (
      .in(par_done_reg21_in),
      .write_en(par_done_reg21_write_en),
      .clk(clk),
      .out(par_done_reg21_out),
      .done(par_done_reg21_done)
  );
  
  std_reg #(1) par_done_reg22 (
      .in(par_done_reg22_in),
      .write_en(par_done_reg22_write_en),
      .clk(clk),
      .out(par_done_reg22_out),
      .done(par_done_reg22_done)
  );
  
  std_reg #(1) par_done_reg23 (
      .in(par_done_reg23_in),
      .write_en(par_done_reg23_write_en),
      .clk(clk),
      .out(par_done_reg23_out),
      .done(par_done_reg23_done)
  );
  
  std_reg #(1) par_done_reg24 (
      .in(par_done_reg24_in),
      .write_en(par_done_reg24_write_en),
      .clk(clk),
      .out(par_done_reg24_out),
      .done(par_done_reg24_done)
  );
  
  std_reg #(1) par_done_reg25 (
      .in(par_done_reg25_in),
      .write_en(par_done_reg25_write_en),
      .clk(clk),
      .out(par_done_reg25_out),
      .done(par_done_reg25_done)
  );
  
  std_reg #(1) par_done_reg26 (
      .in(par_done_reg26_in),
      .write_en(par_done_reg26_write_en),
      .clk(clk),
      .out(par_done_reg26_out),
      .done(par_done_reg26_done)
  );
  
  std_reg #(1) par_reset5 (
      .in(par_reset5_in),
      .write_en(par_reset5_write_en),
      .clk(clk),
      .out(par_reset5_out),
      .done(par_reset5_done)
  );
  
  std_reg #(1) par_done_reg27 (
      .in(par_done_reg27_in),
      .write_en(par_done_reg27_write_en),
      .clk(clk),
      .out(par_done_reg27_out),
      .done(par_done_reg27_done)
  );
  
  std_reg #(1) par_done_reg28 (
      .in(par_done_reg28_in),
      .write_en(par_done_reg28_write_en),
      .clk(clk),
      .out(par_done_reg28_out),
      .done(par_done_reg28_done)
  );
  
  std_reg #(1) par_done_reg29 (
      .in(par_done_reg29_in),
      .write_en(par_done_reg29_write_en),
      .clk(clk),
      .out(par_done_reg29_out),
      .done(par_done_reg29_done)
  );
  
  std_reg #(1) par_done_reg30 (
      .in(par_done_reg30_in),
      .write_en(par_done_reg30_write_en),
      .clk(clk),
      .out(par_done_reg30_out),
      .done(par_done_reg30_done)
  );
  
  std_reg #(1) par_done_reg31 (
      .in(par_done_reg31_in),
      .write_en(par_done_reg31_write_en),
      .clk(clk),
      .out(par_done_reg31_out),
      .done(par_done_reg31_done)
  );
  
  std_reg #(1) par_done_reg32 (
      .in(par_done_reg32_in),
      .write_en(par_done_reg32_write_en),
      .clk(clk),
      .out(par_done_reg32_out),
      .done(par_done_reg32_done)
  );
  
  std_reg #(1) par_done_reg33 (
      .in(par_done_reg33_in),
      .write_en(par_done_reg33_write_en),
      .clk(clk),
      .out(par_done_reg33_out),
      .done(par_done_reg33_done)
  );
  
  std_reg #(1) par_done_reg34 (
      .in(par_done_reg34_in),
      .write_en(par_done_reg34_write_en),
      .clk(clk),
      .out(par_done_reg34_out),
      .done(par_done_reg34_done)
  );
  
  std_reg #(1) par_done_reg35 (
      .in(par_done_reg35_in),
      .write_en(par_done_reg35_write_en),
      .clk(clk),
      .out(par_done_reg35_out),
      .done(par_done_reg35_done)
  );
  
  std_reg #(1) par_reset6 (
      .in(par_reset6_in),
      .write_en(par_reset6_write_en),
      .clk(clk),
      .out(par_reset6_out),
      .done(par_reset6_done)
  );
  
  std_reg #(1) par_done_reg36 (
      .in(par_done_reg36_in),
      .write_en(par_done_reg36_write_en),
      .clk(clk),
      .out(par_done_reg36_out),
      .done(par_done_reg36_done)
  );
  
  std_reg #(1) par_done_reg37 (
      .in(par_done_reg37_in),
      .write_en(par_done_reg37_write_en),
      .clk(clk),
      .out(par_done_reg37_out),
      .done(par_done_reg37_done)
  );
  
  std_reg #(1) par_done_reg38 (
      .in(par_done_reg38_in),
      .write_en(par_done_reg38_write_en),
      .clk(clk),
      .out(par_done_reg38_out),
      .done(par_done_reg38_done)
  );
  
  std_reg #(1) par_done_reg39 (
      .in(par_done_reg39_in),
      .write_en(par_done_reg39_write_en),
      .clk(clk),
      .out(par_done_reg39_out),
      .done(par_done_reg39_done)
  );
  
  std_reg #(1) par_done_reg40 (
      .in(par_done_reg40_in),
      .write_en(par_done_reg40_write_en),
      .clk(clk),
      .out(par_done_reg40_out),
      .done(par_done_reg40_done)
  );
  
  std_reg #(1) par_done_reg41 (
      .in(par_done_reg41_in),
      .write_en(par_done_reg41_write_en),
      .clk(clk),
      .out(par_done_reg41_out),
      .done(par_done_reg41_done)
  );
  
  std_reg #(1) par_done_reg42 (
      .in(par_done_reg42_in),
      .write_en(par_done_reg42_write_en),
      .clk(clk),
      .out(par_done_reg42_out),
      .done(par_done_reg42_done)
  );
  
  std_reg #(1) par_done_reg43 (
      .in(par_done_reg43_in),
      .write_en(par_done_reg43_write_en),
      .clk(clk),
      .out(par_done_reg43_out),
      .done(par_done_reg43_done)
  );
  
  std_reg #(1) par_done_reg44 (
      .in(par_done_reg44_in),
      .write_en(par_done_reg44_write_en),
      .clk(clk),
      .out(par_done_reg44_out),
      .done(par_done_reg44_done)
  );
  
  std_reg #(1) par_done_reg45 (
      .in(par_done_reg45_in),
      .write_en(par_done_reg45_write_en),
      .clk(clk),
      .out(par_done_reg45_out),
      .done(par_done_reg45_done)
  );
  
  std_reg #(1) par_done_reg46 (
      .in(par_done_reg46_in),
      .write_en(par_done_reg46_write_en),
      .clk(clk),
      .out(par_done_reg46_out),
      .done(par_done_reg46_done)
  );
  
  std_reg #(1) par_done_reg47 (
      .in(par_done_reg47_in),
      .write_en(par_done_reg47_write_en),
      .clk(clk),
      .out(par_done_reg47_out),
      .done(par_done_reg47_done)
  );
  
  std_reg #(1) par_reset7 (
      .in(par_reset7_in),
      .write_en(par_reset7_write_en),
      .clk(clk),
      .out(par_reset7_out),
      .done(par_reset7_done)
  );
  
  std_reg #(1) par_done_reg48 (
      .in(par_done_reg48_in),
      .write_en(par_done_reg48_write_en),
      .clk(clk),
      .out(par_done_reg48_out),
      .done(par_done_reg48_done)
  );
  
  std_reg #(1) par_done_reg49 (
      .in(par_done_reg49_in),
      .write_en(par_done_reg49_write_en),
      .clk(clk),
      .out(par_done_reg49_out),
      .done(par_done_reg49_done)
  );
  
  std_reg #(1) par_done_reg50 (
      .in(par_done_reg50_in),
      .write_en(par_done_reg50_write_en),
      .clk(clk),
      .out(par_done_reg50_out),
      .done(par_done_reg50_done)
  );
  
  std_reg #(1) par_done_reg51 (
      .in(par_done_reg51_in),
      .write_en(par_done_reg51_write_en),
      .clk(clk),
      .out(par_done_reg51_out),
      .done(par_done_reg51_done)
  );
  
  std_reg #(1) par_done_reg52 (
      .in(par_done_reg52_in),
      .write_en(par_done_reg52_write_en),
      .clk(clk),
      .out(par_done_reg52_out),
      .done(par_done_reg52_done)
  );
  
  std_reg #(1) par_done_reg53 (
      .in(par_done_reg53_in),
      .write_en(par_done_reg53_write_en),
      .clk(clk),
      .out(par_done_reg53_out),
      .done(par_done_reg53_done)
  );
  
  std_reg #(1) par_done_reg54 (
      .in(par_done_reg54_in),
      .write_en(par_done_reg54_write_en),
      .clk(clk),
      .out(par_done_reg54_out),
      .done(par_done_reg54_done)
  );
  
  std_reg #(1) par_done_reg55 (
      .in(par_done_reg55_in),
      .write_en(par_done_reg55_write_en),
      .clk(clk),
      .out(par_done_reg55_out),
      .done(par_done_reg55_done)
  );
  
  std_reg #(1) par_done_reg56 (
      .in(par_done_reg56_in),
      .write_en(par_done_reg56_write_en),
      .clk(clk),
      .out(par_done_reg56_out),
      .done(par_done_reg56_done)
  );
  
  std_reg #(1) par_done_reg57 (
      .in(par_done_reg57_in),
      .write_en(par_done_reg57_write_en),
      .clk(clk),
      .out(par_done_reg57_out),
      .done(par_done_reg57_done)
  );
  
  std_reg #(1) par_done_reg58 (
      .in(par_done_reg58_in),
      .write_en(par_done_reg58_write_en),
      .clk(clk),
      .out(par_done_reg58_out),
      .done(par_done_reg58_done)
  );
  
  std_reg #(1) par_done_reg59 (
      .in(par_done_reg59_in),
      .write_en(par_done_reg59_write_en),
      .clk(clk),
      .out(par_done_reg59_out),
      .done(par_done_reg59_done)
  );
  
  std_reg #(1) par_done_reg60 (
      .in(par_done_reg60_in),
      .write_en(par_done_reg60_write_en),
      .clk(clk),
      .out(par_done_reg60_out),
      .done(par_done_reg60_done)
  );
  
  std_reg #(1) par_done_reg61 (
      .in(par_done_reg61_in),
      .write_en(par_done_reg61_write_en),
      .clk(clk),
      .out(par_done_reg61_out),
      .done(par_done_reg61_done)
  );
  
  std_reg #(1) par_reset8 (
      .in(par_reset8_in),
      .write_en(par_reset8_write_en),
      .clk(clk),
      .out(par_reset8_out),
      .done(par_reset8_done)
  );
  
  std_reg #(1) par_done_reg62 (
      .in(par_done_reg62_in),
      .write_en(par_done_reg62_write_en),
      .clk(clk),
      .out(par_done_reg62_out),
      .done(par_done_reg62_done)
  );
  
  std_reg #(1) par_done_reg63 (
      .in(par_done_reg63_in),
      .write_en(par_done_reg63_write_en),
      .clk(clk),
      .out(par_done_reg63_out),
      .done(par_done_reg63_done)
  );
  
  std_reg #(1) par_done_reg64 (
      .in(par_done_reg64_in),
      .write_en(par_done_reg64_write_en),
      .clk(clk),
      .out(par_done_reg64_out),
      .done(par_done_reg64_done)
  );
  
  std_reg #(1) par_done_reg65 (
      .in(par_done_reg65_in),
      .write_en(par_done_reg65_write_en),
      .clk(clk),
      .out(par_done_reg65_out),
      .done(par_done_reg65_done)
  );
  
  std_reg #(1) par_done_reg66 (
      .in(par_done_reg66_in),
      .write_en(par_done_reg66_write_en),
      .clk(clk),
      .out(par_done_reg66_out),
      .done(par_done_reg66_done)
  );
  
  std_reg #(1) par_done_reg67 (
      .in(par_done_reg67_in),
      .write_en(par_done_reg67_write_en),
      .clk(clk),
      .out(par_done_reg67_out),
      .done(par_done_reg67_done)
  );
  
  std_reg #(1) par_done_reg68 (
      .in(par_done_reg68_in),
      .write_en(par_done_reg68_write_en),
      .clk(clk),
      .out(par_done_reg68_out),
      .done(par_done_reg68_done)
  );
  
  std_reg #(1) par_done_reg69 (
      .in(par_done_reg69_in),
      .write_en(par_done_reg69_write_en),
      .clk(clk),
      .out(par_done_reg69_out),
      .done(par_done_reg69_done)
  );
  
  std_reg #(1) par_done_reg70 (
      .in(par_done_reg70_in),
      .write_en(par_done_reg70_write_en),
      .clk(clk),
      .out(par_done_reg70_out),
      .done(par_done_reg70_done)
  );
  
  std_reg #(1) par_done_reg71 (
      .in(par_done_reg71_in),
      .write_en(par_done_reg71_write_en),
      .clk(clk),
      .out(par_done_reg71_out),
      .done(par_done_reg71_done)
  );
  
  std_reg #(1) par_done_reg72 (
      .in(par_done_reg72_in),
      .write_en(par_done_reg72_write_en),
      .clk(clk),
      .out(par_done_reg72_out),
      .done(par_done_reg72_done)
  );
  
  std_reg #(1) par_done_reg73 (
      .in(par_done_reg73_in),
      .write_en(par_done_reg73_write_en),
      .clk(clk),
      .out(par_done_reg73_out),
      .done(par_done_reg73_done)
  );
  
  std_reg #(1) par_done_reg74 (
      .in(par_done_reg74_in),
      .write_en(par_done_reg74_write_en),
      .clk(clk),
      .out(par_done_reg74_out),
      .done(par_done_reg74_done)
  );
  
  std_reg #(1) par_done_reg75 (
      .in(par_done_reg75_in),
      .write_en(par_done_reg75_write_en),
      .clk(clk),
      .out(par_done_reg75_out),
      .done(par_done_reg75_done)
  );
  
  std_reg #(1) par_done_reg76 (
      .in(par_done_reg76_in),
      .write_en(par_done_reg76_write_en),
      .clk(clk),
      .out(par_done_reg76_out),
      .done(par_done_reg76_done)
  );
  
  std_reg #(1) par_done_reg77 (
      .in(par_done_reg77_in),
      .write_en(par_done_reg77_write_en),
      .clk(clk),
      .out(par_done_reg77_out),
      .done(par_done_reg77_done)
  );
  
  std_reg #(1) par_done_reg78 (
      .in(par_done_reg78_in),
      .write_en(par_done_reg78_write_en),
      .clk(clk),
      .out(par_done_reg78_out),
      .done(par_done_reg78_done)
  );
  
  std_reg #(1) par_done_reg79 (
      .in(par_done_reg79_in),
      .write_en(par_done_reg79_write_en),
      .clk(clk),
      .out(par_done_reg79_out),
      .done(par_done_reg79_done)
  );
  
  std_reg #(1) par_done_reg80 (
      .in(par_done_reg80_in),
      .write_en(par_done_reg80_write_en),
      .clk(clk),
      .out(par_done_reg80_out),
      .done(par_done_reg80_done)
  );
  
  std_reg #(1) par_done_reg81 (
      .in(par_done_reg81_in),
      .write_en(par_done_reg81_write_en),
      .clk(clk),
      .out(par_done_reg81_out),
      .done(par_done_reg81_done)
  );
  
  std_reg #(1) par_reset9 (
      .in(par_reset9_in),
      .write_en(par_reset9_write_en),
      .clk(clk),
      .out(par_reset9_out),
      .done(par_reset9_done)
  );
  
  std_reg #(1) par_done_reg82 (
      .in(par_done_reg82_in),
      .write_en(par_done_reg82_write_en),
      .clk(clk),
      .out(par_done_reg82_out),
      .done(par_done_reg82_done)
  );
  
  std_reg #(1) par_done_reg83 (
      .in(par_done_reg83_in),
      .write_en(par_done_reg83_write_en),
      .clk(clk),
      .out(par_done_reg83_out),
      .done(par_done_reg83_done)
  );
  
  std_reg #(1) par_done_reg84 (
      .in(par_done_reg84_in),
      .write_en(par_done_reg84_write_en),
      .clk(clk),
      .out(par_done_reg84_out),
      .done(par_done_reg84_done)
  );
  
  std_reg #(1) par_done_reg85 (
      .in(par_done_reg85_in),
      .write_en(par_done_reg85_write_en),
      .clk(clk),
      .out(par_done_reg85_out),
      .done(par_done_reg85_done)
  );
  
  std_reg #(1) par_done_reg86 (
      .in(par_done_reg86_in),
      .write_en(par_done_reg86_write_en),
      .clk(clk),
      .out(par_done_reg86_out),
      .done(par_done_reg86_done)
  );
  
  std_reg #(1) par_done_reg87 (
      .in(par_done_reg87_in),
      .write_en(par_done_reg87_write_en),
      .clk(clk),
      .out(par_done_reg87_out),
      .done(par_done_reg87_done)
  );
  
  std_reg #(1) par_done_reg88 (
      .in(par_done_reg88_in),
      .write_en(par_done_reg88_write_en),
      .clk(clk),
      .out(par_done_reg88_out),
      .done(par_done_reg88_done)
  );
  
  std_reg #(1) par_done_reg89 (
      .in(par_done_reg89_in),
      .write_en(par_done_reg89_write_en),
      .clk(clk),
      .out(par_done_reg89_out),
      .done(par_done_reg89_done)
  );
  
  std_reg #(1) par_done_reg90 (
      .in(par_done_reg90_in),
      .write_en(par_done_reg90_write_en),
      .clk(clk),
      .out(par_done_reg90_out),
      .done(par_done_reg90_done)
  );
  
  std_reg #(1) par_done_reg91 (
      .in(par_done_reg91_in),
      .write_en(par_done_reg91_write_en),
      .clk(clk),
      .out(par_done_reg91_out),
      .done(par_done_reg91_done)
  );
  
  std_reg #(1) par_done_reg92 (
      .in(par_done_reg92_in),
      .write_en(par_done_reg92_write_en),
      .clk(clk),
      .out(par_done_reg92_out),
      .done(par_done_reg92_done)
  );
  
  std_reg #(1) par_done_reg93 (
      .in(par_done_reg93_in),
      .write_en(par_done_reg93_write_en),
      .clk(clk),
      .out(par_done_reg93_out),
      .done(par_done_reg93_done)
  );
  
  std_reg #(1) par_done_reg94 (
      .in(par_done_reg94_in),
      .write_en(par_done_reg94_write_en),
      .clk(clk),
      .out(par_done_reg94_out),
      .done(par_done_reg94_done)
  );
  
  std_reg #(1) par_done_reg95 (
      .in(par_done_reg95_in),
      .write_en(par_done_reg95_write_en),
      .clk(clk),
      .out(par_done_reg95_out),
      .done(par_done_reg95_done)
  );
  
  std_reg #(1) par_done_reg96 (
      .in(par_done_reg96_in),
      .write_en(par_done_reg96_write_en),
      .clk(clk),
      .out(par_done_reg96_out),
      .done(par_done_reg96_done)
  );
  
  std_reg #(1) par_done_reg97 (
      .in(par_done_reg97_in),
      .write_en(par_done_reg97_write_en),
      .clk(clk),
      .out(par_done_reg97_out),
      .done(par_done_reg97_done)
  );
  
  std_reg #(1) par_done_reg98 (
      .in(par_done_reg98_in),
      .write_en(par_done_reg98_write_en),
      .clk(clk),
      .out(par_done_reg98_out),
      .done(par_done_reg98_done)
  );
  
  std_reg #(1) par_done_reg99 (
      .in(par_done_reg99_in),
      .write_en(par_done_reg99_write_en),
      .clk(clk),
      .out(par_done_reg99_out),
      .done(par_done_reg99_done)
  );
  
  std_reg #(1) par_done_reg100 (
      .in(par_done_reg100_in),
      .write_en(par_done_reg100_write_en),
      .clk(clk),
      .out(par_done_reg100_out),
      .done(par_done_reg100_done)
  );
  
  std_reg #(1) par_done_reg101 (
      .in(par_done_reg101_in),
      .write_en(par_done_reg101_write_en),
      .clk(clk),
      .out(par_done_reg101_out),
      .done(par_done_reg101_done)
  );
  
  std_reg #(1) par_reset10 (
      .in(par_reset10_in),
      .write_en(par_reset10_write_en),
      .clk(clk),
      .out(par_reset10_out),
      .done(par_reset10_done)
  );
  
  std_reg #(1) par_done_reg102 (
      .in(par_done_reg102_in),
      .write_en(par_done_reg102_write_en),
      .clk(clk),
      .out(par_done_reg102_out),
      .done(par_done_reg102_done)
  );
  
  std_reg #(1) par_done_reg103 (
      .in(par_done_reg103_in),
      .write_en(par_done_reg103_write_en),
      .clk(clk),
      .out(par_done_reg103_out),
      .done(par_done_reg103_done)
  );
  
  std_reg #(1) par_done_reg104 (
      .in(par_done_reg104_in),
      .write_en(par_done_reg104_write_en),
      .clk(clk),
      .out(par_done_reg104_out),
      .done(par_done_reg104_done)
  );
  
  std_reg #(1) par_done_reg105 (
      .in(par_done_reg105_in),
      .write_en(par_done_reg105_write_en),
      .clk(clk),
      .out(par_done_reg105_out),
      .done(par_done_reg105_done)
  );
  
  std_reg #(1) par_done_reg106 (
      .in(par_done_reg106_in),
      .write_en(par_done_reg106_write_en),
      .clk(clk),
      .out(par_done_reg106_out),
      .done(par_done_reg106_done)
  );
  
  std_reg #(1) par_done_reg107 (
      .in(par_done_reg107_in),
      .write_en(par_done_reg107_write_en),
      .clk(clk),
      .out(par_done_reg107_out),
      .done(par_done_reg107_done)
  );
  
  std_reg #(1) par_done_reg108 (
      .in(par_done_reg108_in),
      .write_en(par_done_reg108_write_en),
      .clk(clk),
      .out(par_done_reg108_out),
      .done(par_done_reg108_done)
  );
  
  std_reg #(1) par_done_reg109 (
      .in(par_done_reg109_in),
      .write_en(par_done_reg109_write_en),
      .clk(clk),
      .out(par_done_reg109_out),
      .done(par_done_reg109_done)
  );
  
  std_reg #(1) par_done_reg110 (
      .in(par_done_reg110_in),
      .write_en(par_done_reg110_write_en),
      .clk(clk),
      .out(par_done_reg110_out),
      .done(par_done_reg110_done)
  );
  
  std_reg #(1) par_done_reg111 (
      .in(par_done_reg111_in),
      .write_en(par_done_reg111_write_en),
      .clk(clk),
      .out(par_done_reg111_out),
      .done(par_done_reg111_done)
  );
  
  std_reg #(1) par_done_reg112 (
      .in(par_done_reg112_in),
      .write_en(par_done_reg112_write_en),
      .clk(clk),
      .out(par_done_reg112_out),
      .done(par_done_reg112_done)
  );
  
  std_reg #(1) par_done_reg113 (
      .in(par_done_reg113_in),
      .write_en(par_done_reg113_write_en),
      .clk(clk),
      .out(par_done_reg113_out),
      .done(par_done_reg113_done)
  );
  
  std_reg #(1) par_done_reg114 (
      .in(par_done_reg114_in),
      .write_en(par_done_reg114_write_en),
      .clk(clk),
      .out(par_done_reg114_out),
      .done(par_done_reg114_done)
  );
  
  std_reg #(1) par_done_reg115 (
      .in(par_done_reg115_in),
      .write_en(par_done_reg115_write_en),
      .clk(clk),
      .out(par_done_reg115_out),
      .done(par_done_reg115_done)
  );
  
  std_reg #(1) par_done_reg116 (
      .in(par_done_reg116_in),
      .write_en(par_done_reg116_write_en),
      .clk(clk),
      .out(par_done_reg116_out),
      .done(par_done_reg116_done)
  );
  
  std_reg #(1) par_done_reg117 (
      .in(par_done_reg117_in),
      .write_en(par_done_reg117_write_en),
      .clk(clk),
      .out(par_done_reg117_out),
      .done(par_done_reg117_done)
  );
  
  std_reg #(1) par_done_reg118 (
      .in(par_done_reg118_in),
      .write_en(par_done_reg118_write_en),
      .clk(clk),
      .out(par_done_reg118_out),
      .done(par_done_reg118_done)
  );
  
  std_reg #(1) par_done_reg119 (
      .in(par_done_reg119_in),
      .write_en(par_done_reg119_write_en),
      .clk(clk),
      .out(par_done_reg119_out),
      .done(par_done_reg119_done)
  );
  
  std_reg #(1) par_done_reg120 (
      .in(par_done_reg120_in),
      .write_en(par_done_reg120_write_en),
      .clk(clk),
      .out(par_done_reg120_out),
      .done(par_done_reg120_done)
  );
  
  std_reg #(1) par_done_reg121 (
      .in(par_done_reg121_in),
      .write_en(par_done_reg121_write_en),
      .clk(clk),
      .out(par_done_reg121_out),
      .done(par_done_reg121_done)
  );
  
  std_reg #(1) par_done_reg122 (
      .in(par_done_reg122_in),
      .write_en(par_done_reg122_write_en),
      .clk(clk),
      .out(par_done_reg122_out),
      .done(par_done_reg122_done)
  );
  
  std_reg #(1) par_done_reg123 (
      .in(par_done_reg123_in),
      .write_en(par_done_reg123_write_en),
      .clk(clk),
      .out(par_done_reg123_out),
      .done(par_done_reg123_done)
  );
  
  std_reg #(1) par_done_reg124 (
      .in(par_done_reg124_in),
      .write_en(par_done_reg124_write_en),
      .clk(clk),
      .out(par_done_reg124_out),
      .done(par_done_reg124_done)
  );
  
  std_reg #(1) par_done_reg125 (
      .in(par_done_reg125_in),
      .write_en(par_done_reg125_write_en),
      .clk(clk),
      .out(par_done_reg125_out),
      .done(par_done_reg125_done)
  );
  
  std_reg #(1) par_done_reg126 (
      .in(par_done_reg126_in),
      .write_en(par_done_reg126_write_en),
      .clk(clk),
      .out(par_done_reg126_out),
      .done(par_done_reg126_done)
  );
  
  std_reg #(1) par_done_reg127 (
      .in(par_done_reg127_in),
      .write_en(par_done_reg127_write_en),
      .clk(clk),
      .out(par_done_reg127_out),
      .done(par_done_reg127_done)
  );
  
  std_reg #(1) par_done_reg128 (
      .in(par_done_reg128_in),
      .write_en(par_done_reg128_write_en),
      .clk(clk),
      .out(par_done_reg128_out),
      .done(par_done_reg128_done)
  );
  
  std_reg #(1) par_done_reg129 (
      .in(par_done_reg129_in),
      .write_en(par_done_reg129_write_en),
      .clk(clk),
      .out(par_done_reg129_out),
      .done(par_done_reg129_done)
  );
  
  std_reg #(1) par_done_reg130 (
      .in(par_done_reg130_in),
      .write_en(par_done_reg130_write_en),
      .clk(clk),
      .out(par_done_reg130_out),
      .done(par_done_reg130_done)
  );
  
  std_reg #(1) par_done_reg131 (
      .in(par_done_reg131_in),
      .write_en(par_done_reg131_write_en),
      .clk(clk),
      .out(par_done_reg131_out),
      .done(par_done_reg131_done)
  );
  
  std_reg #(1) par_reset11 (
      .in(par_reset11_in),
      .write_en(par_reset11_write_en),
      .clk(clk),
      .out(par_reset11_out),
      .done(par_reset11_done)
  );
  
  std_reg #(1) par_done_reg132 (
      .in(par_done_reg132_in),
      .write_en(par_done_reg132_write_en),
      .clk(clk),
      .out(par_done_reg132_out),
      .done(par_done_reg132_done)
  );
  
  std_reg #(1) par_done_reg133 (
      .in(par_done_reg133_in),
      .write_en(par_done_reg133_write_en),
      .clk(clk),
      .out(par_done_reg133_out),
      .done(par_done_reg133_done)
  );
  
  std_reg #(1) par_done_reg134 (
      .in(par_done_reg134_in),
      .write_en(par_done_reg134_write_en),
      .clk(clk),
      .out(par_done_reg134_out),
      .done(par_done_reg134_done)
  );
  
  std_reg #(1) par_done_reg135 (
      .in(par_done_reg135_in),
      .write_en(par_done_reg135_write_en),
      .clk(clk),
      .out(par_done_reg135_out),
      .done(par_done_reg135_done)
  );
  
  std_reg #(1) par_done_reg136 (
      .in(par_done_reg136_in),
      .write_en(par_done_reg136_write_en),
      .clk(clk),
      .out(par_done_reg136_out),
      .done(par_done_reg136_done)
  );
  
  std_reg #(1) par_done_reg137 (
      .in(par_done_reg137_in),
      .write_en(par_done_reg137_write_en),
      .clk(clk),
      .out(par_done_reg137_out),
      .done(par_done_reg137_done)
  );
  
  std_reg #(1) par_done_reg138 (
      .in(par_done_reg138_in),
      .write_en(par_done_reg138_write_en),
      .clk(clk),
      .out(par_done_reg138_out),
      .done(par_done_reg138_done)
  );
  
  std_reg #(1) par_done_reg139 (
      .in(par_done_reg139_in),
      .write_en(par_done_reg139_write_en),
      .clk(clk),
      .out(par_done_reg139_out),
      .done(par_done_reg139_done)
  );
  
  std_reg #(1) par_done_reg140 (
      .in(par_done_reg140_in),
      .write_en(par_done_reg140_write_en),
      .clk(clk),
      .out(par_done_reg140_out),
      .done(par_done_reg140_done)
  );
  
  std_reg #(1) par_done_reg141 (
      .in(par_done_reg141_in),
      .write_en(par_done_reg141_write_en),
      .clk(clk),
      .out(par_done_reg141_out),
      .done(par_done_reg141_done)
  );
  
  std_reg #(1) par_done_reg142 (
      .in(par_done_reg142_in),
      .write_en(par_done_reg142_write_en),
      .clk(clk),
      .out(par_done_reg142_out),
      .done(par_done_reg142_done)
  );
  
  std_reg #(1) par_done_reg143 (
      .in(par_done_reg143_in),
      .write_en(par_done_reg143_write_en),
      .clk(clk),
      .out(par_done_reg143_out),
      .done(par_done_reg143_done)
  );
  
  std_reg #(1) par_done_reg144 (
      .in(par_done_reg144_in),
      .write_en(par_done_reg144_write_en),
      .clk(clk),
      .out(par_done_reg144_out),
      .done(par_done_reg144_done)
  );
  
  std_reg #(1) par_done_reg145 (
      .in(par_done_reg145_in),
      .write_en(par_done_reg145_write_en),
      .clk(clk),
      .out(par_done_reg145_out),
      .done(par_done_reg145_done)
  );
  
  std_reg #(1) par_done_reg146 (
      .in(par_done_reg146_in),
      .write_en(par_done_reg146_write_en),
      .clk(clk),
      .out(par_done_reg146_out),
      .done(par_done_reg146_done)
  );
  
  std_reg #(1) par_done_reg147 (
      .in(par_done_reg147_in),
      .write_en(par_done_reg147_write_en),
      .clk(clk),
      .out(par_done_reg147_out),
      .done(par_done_reg147_done)
  );
  
  std_reg #(1) par_done_reg148 (
      .in(par_done_reg148_in),
      .write_en(par_done_reg148_write_en),
      .clk(clk),
      .out(par_done_reg148_out),
      .done(par_done_reg148_done)
  );
  
  std_reg #(1) par_done_reg149 (
      .in(par_done_reg149_in),
      .write_en(par_done_reg149_write_en),
      .clk(clk),
      .out(par_done_reg149_out),
      .done(par_done_reg149_done)
  );
  
  std_reg #(1) par_done_reg150 (
      .in(par_done_reg150_in),
      .write_en(par_done_reg150_write_en),
      .clk(clk),
      .out(par_done_reg150_out),
      .done(par_done_reg150_done)
  );
  
  std_reg #(1) par_done_reg151 (
      .in(par_done_reg151_in),
      .write_en(par_done_reg151_write_en),
      .clk(clk),
      .out(par_done_reg151_out),
      .done(par_done_reg151_done)
  );
  
  std_reg #(1) par_done_reg152 (
      .in(par_done_reg152_in),
      .write_en(par_done_reg152_write_en),
      .clk(clk),
      .out(par_done_reg152_out),
      .done(par_done_reg152_done)
  );
  
  std_reg #(1) par_done_reg153 (
      .in(par_done_reg153_in),
      .write_en(par_done_reg153_write_en),
      .clk(clk),
      .out(par_done_reg153_out),
      .done(par_done_reg153_done)
  );
  
  std_reg #(1) par_done_reg154 (
      .in(par_done_reg154_in),
      .write_en(par_done_reg154_write_en),
      .clk(clk),
      .out(par_done_reg154_out),
      .done(par_done_reg154_done)
  );
  
  std_reg #(1) par_done_reg155 (
      .in(par_done_reg155_in),
      .write_en(par_done_reg155_write_en),
      .clk(clk),
      .out(par_done_reg155_out),
      .done(par_done_reg155_done)
  );
  
  std_reg #(1) par_done_reg156 (
      .in(par_done_reg156_in),
      .write_en(par_done_reg156_write_en),
      .clk(clk),
      .out(par_done_reg156_out),
      .done(par_done_reg156_done)
  );
  
  std_reg #(1) par_done_reg157 (
      .in(par_done_reg157_in),
      .write_en(par_done_reg157_write_en),
      .clk(clk),
      .out(par_done_reg157_out),
      .done(par_done_reg157_done)
  );
  
  std_reg #(1) par_done_reg158 (
      .in(par_done_reg158_in),
      .write_en(par_done_reg158_write_en),
      .clk(clk),
      .out(par_done_reg158_out),
      .done(par_done_reg158_done)
  );
  
  std_reg #(1) par_reset12 (
      .in(par_reset12_in),
      .write_en(par_reset12_write_en),
      .clk(clk),
      .out(par_reset12_out),
      .done(par_reset12_done)
  );
  
  std_reg #(1) par_done_reg159 (
      .in(par_done_reg159_in),
      .write_en(par_done_reg159_write_en),
      .clk(clk),
      .out(par_done_reg159_out),
      .done(par_done_reg159_done)
  );
  
  std_reg #(1) par_done_reg160 (
      .in(par_done_reg160_in),
      .write_en(par_done_reg160_write_en),
      .clk(clk),
      .out(par_done_reg160_out),
      .done(par_done_reg160_done)
  );
  
  std_reg #(1) par_done_reg161 (
      .in(par_done_reg161_in),
      .write_en(par_done_reg161_write_en),
      .clk(clk),
      .out(par_done_reg161_out),
      .done(par_done_reg161_done)
  );
  
  std_reg #(1) par_done_reg162 (
      .in(par_done_reg162_in),
      .write_en(par_done_reg162_write_en),
      .clk(clk),
      .out(par_done_reg162_out),
      .done(par_done_reg162_done)
  );
  
  std_reg #(1) par_done_reg163 (
      .in(par_done_reg163_in),
      .write_en(par_done_reg163_write_en),
      .clk(clk),
      .out(par_done_reg163_out),
      .done(par_done_reg163_done)
  );
  
  std_reg #(1) par_done_reg164 (
      .in(par_done_reg164_in),
      .write_en(par_done_reg164_write_en),
      .clk(clk),
      .out(par_done_reg164_out),
      .done(par_done_reg164_done)
  );
  
  std_reg #(1) par_done_reg165 (
      .in(par_done_reg165_in),
      .write_en(par_done_reg165_write_en),
      .clk(clk),
      .out(par_done_reg165_out),
      .done(par_done_reg165_done)
  );
  
  std_reg #(1) par_done_reg166 (
      .in(par_done_reg166_in),
      .write_en(par_done_reg166_write_en),
      .clk(clk),
      .out(par_done_reg166_out),
      .done(par_done_reg166_done)
  );
  
  std_reg #(1) par_done_reg167 (
      .in(par_done_reg167_in),
      .write_en(par_done_reg167_write_en),
      .clk(clk),
      .out(par_done_reg167_out),
      .done(par_done_reg167_done)
  );
  
  std_reg #(1) par_done_reg168 (
      .in(par_done_reg168_in),
      .write_en(par_done_reg168_write_en),
      .clk(clk),
      .out(par_done_reg168_out),
      .done(par_done_reg168_done)
  );
  
  std_reg #(1) par_done_reg169 (
      .in(par_done_reg169_in),
      .write_en(par_done_reg169_write_en),
      .clk(clk),
      .out(par_done_reg169_out),
      .done(par_done_reg169_done)
  );
  
  std_reg #(1) par_done_reg170 (
      .in(par_done_reg170_in),
      .write_en(par_done_reg170_write_en),
      .clk(clk),
      .out(par_done_reg170_out),
      .done(par_done_reg170_done)
  );
  
  std_reg #(1) par_done_reg171 (
      .in(par_done_reg171_in),
      .write_en(par_done_reg171_write_en),
      .clk(clk),
      .out(par_done_reg171_out),
      .done(par_done_reg171_done)
  );
  
  std_reg #(1) par_done_reg172 (
      .in(par_done_reg172_in),
      .write_en(par_done_reg172_write_en),
      .clk(clk),
      .out(par_done_reg172_out),
      .done(par_done_reg172_done)
  );
  
  std_reg #(1) par_done_reg173 (
      .in(par_done_reg173_in),
      .write_en(par_done_reg173_write_en),
      .clk(clk),
      .out(par_done_reg173_out),
      .done(par_done_reg173_done)
  );
  
  std_reg #(1) par_done_reg174 (
      .in(par_done_reg174_in),
      .write_en(par_done_reg174_write_en),
      .clk(clk),
      .out(par_done_reg174_out),
      .done(par_done_reg174_done)
  );
  
  std_reg #(1) par_done_reg175 (
      .in(par_done_reg175_in),
      .write_en(par_done_reg175_write_en),
      .clk(clk),
      .out(par_done_reg175_out),
      .done(par_done_reg175_done)
  );
  
  std_reg #(1) par_done_reg176 (
      .in(par_done_reg176_in),
      .write_en(par_done_reg176_write_en),
      .clk(clk),
      .out(par_done_reg176_out),
      .done(par_done_reg176_done)
  );
  
  std_reg #(1) par_done_reg177 (
      .in(par_done_reg177_in),
      .write_en(par_done_reg177_write_en),
      .clk(clk),
      .out(par_done_reg177_out),
      .done(par_done_reg177_done)
  );
  
  std_reg #(1) par_done_reg178 (
      .in(par_done_reg178_in),
      .write_en(par_done_reg178_write_en),
      .clk(clk),
      .out(par_done_reg178_out),
      .done(par_done_reg178_done)
  );
  
  std_reg #(1) par_done_reg179 (
      .in(par_done_reg179_in),
      .write_en(par_done_reg179_write_en),
      .clk(clk),
      .out(par_done_reg179_out),
      .done(par_done_reg179_done)
  );
  
  std_reg #(1) par_done_reg180 (
      .in(par_done_reg180_in),
      .write_en(par_done_reg180_write_en),
      .clk(clk),
      .out(par_done_reg180_out),
      .done(par_done_reg180_done)
  );
  
  std_reg #(1) par_done_reg181 (
      .in(par_done_reg181_in),
      .write_en(par_done_reg181_write_en),
      .clk(clk),
      .out(par_done_reg181_out),
      .done(par_done_reg181_done)
  );
  
  std_reg #(1) par_done_reg182 (
      .in(par_done_reg182_in),
      .write_en(par_done_reg182_write_en),
      .clk(clk),
      .out(par_done_reg182_out),
      .done(par_done_reg182_done)
  );
  
  std_reg #(1) par_done_reg183 (
      .in(par_done_reg183_in),
      .write_en(par_done_reg183_write_en),
      .clk(clk),
      .out(par_done_reg183_out),
      .done(par_done_reg183_done)
  );
  
  std_reg #(1) par_done_reg184 (
      .in(par_done_reg184_in),
      .write_en(par_done_reg184_write_en),
      .clk(clk),
      .out(par_done_reg184_out),
      .done(par_done_reg184_done)
  );
  
  std_reg #(1) par_done_reg185 (
      .in(par_done_reg185_in),
      .write_en(par_done_reg185_write_en),
      .clk(clk),
      .out(par_done_reg185_out),
      .done(par_done_reg185_done)
  );
  
  std_reg #(1) par_done_reg186 (
      .in(par_done_reg186_in),
      .write_en(par_done_reg186_write_en),
      .clk(clk),
      .out(par_done_reg186_out),
      .done(par_done_reg186_done)
  );
  
  std_reg #(1) par_done_reg187 (
      .in(par_done_reg187_in),
      .write_en(par_done_reg187_write_en),
      .clk(clk),
      .out(par_done_reg187_out),
      .done(par_done_reg187_done)
  );
  
  std_reg #(1) par_done_reg188 (
      .in(par_done_reg188_in),
      .write_en(par_done_reg188_write_en),
      .clk(clk),
      .out(par_done_reg188_out),
      .done(par_done_reg188_done)
  );
  
  std_reg #(1) par_done_reg189 (
      .in(par_done_reg189_in),
      .write_en(par_done_reg189_write_en),
      .clk(clk),
      .out(par_done_reg189_out),
      .done(par_done_reg189_done)
  );
  
  std_reg #(1) par_done_reg190 (
      .in(par_done_reg190_in),
      .write_en(par_done_reg190_write_en),
      .clk(clk),
      .out(par_done_reg190_out),
      .done(par_done_reg190_done)
  );
  
  std_reg #(1) par_done_reg191 (
      .in(par_done_reg191_in),
      .write_en(par_done_reg191_write_en),
      .clk(clk),
      .out(par_done_reg191_out),
      .done(par_done_reg191_done)
  );
  
  std_reg #(1) par_done_reg192 (
      .in(par_done_reg192_in),
      .write_en(par_done_reg192_write_en),
      .clk(clk),
      .out(par_done_reg192_out),
      .done(par_done_reg192_done)
  );
  
  std_reg #(1) par_done_reg193 (
      .in(par_done_reg193_in),
      .write_en(par_done_reg193_write_en),
      .clk(clk),
      .out(par_done_reg193_out),
      .done(par_done_reg193_done)
  );
  
  std_reg #(1) par_done_reg194 (
      .in(par_done_reg194_in),
      .write_en(par_done_reg194_write_en),
      .clk(clk),
      .out(par_done_reg194_out),
      .done(par_done_reg194_done)
  );
  
  std_reg #(1) par_done_reg195 (
      .in(par_done_reg195_in),
      .write_en(par_done_reg195_write_en),
      .clk(clk),
      .out(par_done_reg195_out),
      .done(par_done_reg195_done)
  );
  
  std_reg #(1) par_done_reg196 (
      .in(par_done_reg196_in),
      .write_en(par_done_reg196_write_en),
      .clk(clk),
      .out(par_done_reg196_out),
      .done(par_done_reg196_done)
  );
  
  std_reg #(1) par_done_reg197 (
      .in(par_done_reg197_in),
      .write_en(par_done_reg197_write_en),
      .clk(clk),
      .out(par_done_reg197_out),
      .done(par_done_reg197_done)
  );
  
  std_reg #(1) par_done_reg198 (
      .in(par_done_reg198_in),
      .write_en(par_done_reg198_write_en),
      .clk(clk),
      .out(par_done_reg198_out),
      .done(par_done_reg198_done)
  );
  
  std_reg #(1) par_done_reg199 (
      .in(par_done_reg199_in),
      .write_en(par_done_reg199_write_en),
      .clk(clk),
      .out(par_done_reg199_out),
      .done(par_done_reg199_done)
  );
  
  std_reg #(1) par_done_reg200 (
      .in(par_done_reg200_in),
      .write_en(par_done_reg200_write_en),
      .clk(clk),
      .out(par_done_reg200_out),
      .done(par_done_reg200_done)
  );
  
  std_reg #(1) par_reset13 (
      .in(par_reset13_in),
      .write_en(par_reset13_write_en),
      .clk(clk),
      .out(par_reset13_out),
      .done(par_reset13_done)
  );
  
  std_reg #(1) par_done_reg201 (
      .in(par_done_reg201_in),
      .write_en(par_done_reg201_write_en),
      .clk(clk),
      .out(par_done_reg201_out),
      .done(par_done_reg201_done)
  );
  
  std_reg #(1) par_done_reg202 (
      .in(par_done_reg202_in),
      .write_en(par_done_reg202_write_en),
      .clk(clk),
      .out(par_done_reg202_out),
      .done(par_done_reg202_done)
  );
  
  std_reg #(1) par_done_reg203 (
      .in(par_done_reg203_in),
      .write_en(par_done_reg203_write_en),
      .clk(clk),
      .out(par_done_reg203_out),
      .done(par_done_reg203_done)
  );
  
  std_reg #(1) par_done_reg204 (
      .in(par_done_reg204_in),
      .write_en(par_done_reg204_write_en),
      .clk(clk),
      .out(par_done_reg204_out),
      .done(par_done_reg204_done)
  );
  
  std_reg #(1) par_done_reg205 (
      .in(par_done_reg205_in),
      .write_en(par_done_reg205_write_en),
      .clk(clk),
      .out(par_done_reg205_out),
      .done(par_done_reg205_done)
  );
  
  std_reg #(1) par_done_reg206 (
      .in(par_done_reg206_in),
      .write_en(par_done_reg206_write_en),
      .clk(clk),
      .out(par_done_reg206_out),
      .done(par_done_reg206_done)
  );
  
  std_reg #(1) par_done_reg207 (
      .in(par_done_reg207_in),
      .write_en(par_done_reg207_write_en),
      .clk(clk),
      .out(par_done_reg207_out),
      .done(par_done_reg207_done)
  );
  
  std_reg #(1) par_done_reg208 (
      .in(par_done_reg208_in),
      .write_en(par_done_reg208_write_en),
      .clk(clk),
      .out(par_done_reg208_out),
      .done(par_done_reg208_done)
  );
  
  std_reg #(1) par_done_reg209 (
      .in(par_done_reg209_in),
      .write_en(par_done_reg209_write_en),
      .clk(clk),
      .out(par_done_reg209_out),
      .done(par_done_reg209_done)
  );
  
  std_reg #(1) par_done_reg210 (
      .in(par_done_reg210_in),
      .write_en(par_done_reg210_write_en),
      .clk(clk),
      .out(par_done_reg210_out),
      .done(par_done_reg210_done)
  );
  
  std_reg #(1) par_done_reg211 (
      .in(par_done_reg211_in),
      .write_en(par_done_reg211_write_en),
      .clk(clk),
      .out(par_done_reg211_out),
      .done(par_done_reg211_done)
  );
  
  std_reg #(1) par_done_reg212 (
      .in(par_done_reg212_in),
      .write_en(par_done_reg212_write_en),
      .clk(clk),
      .out(par_done_reg212_out),
      .done(par_done_reg212_done)
  );
  
  std_reg #(1) par_done_reg213 (
      .in(par_done_reg213_in),
      .write_en(par_done_reg213_write_en),
      .clk(clk),
      .out(par_done_reg213_out),
      .done(par_done_reg213_done)
  );
  
  std_reg #(1) par_done_reg214 (
      .in(par_done_reg214_in),
      .write_en(par_done_reg214_write_en),
      .clk(clk),
      .out(par_done_reg214_out),
      .done(par_done_reg214_done)
  );
  
  std_reg #(1) par_done_reg215 (
      .in(par_done_reg215_in),
      .write_en(par_done_reg215_write_en),
      .clk(clk),
      .out(par_done_reg215_out),
      .done(par_done_reg215_done)
  );
  
  std_reg #(1) par_done_reg216 (
      .in(par_done_reg216_in),
      .write_en(par_done_reg216_write_en),
      .clk(clk),
      .out(par_done_reg216_out),
      .done(par_done_reg216_done)
  );
  
  std_reg #(1) par_done_reg217 (
      .in(par_done_reg217_in),
      .write_en(par_done_reg217_write_en),
      .clk(clk),
      .out(par_done_reg217_out),
      .done(par_done_reg217_done)
  );
  
  std_reg #(1) par_done_reg218 (
      .in(par_done_reg218_in),
      .write_en(par_done_reg218_write_en),
      .clk(clk),
      .out(par_done_reg218_out),
      .done(par_done_reg218_done)
  );
  
  std_reg #(1) par_done_reg219 (
      .in(par_done_reg219_in),
      .write_en(par_done_reg219_write_en),
      .clk(clk),
      .out(par_done_reg219_out),
      .done(par_done_reg219_done)
  );
  
  std_reg #(1) par_done_reg220 (
      .in(par_done_reg220_in),
      .write_en(par_done_reg220_write_en),
      .clk(clk),
      .out(par_done_reg220_out),
      .done(par_done_reg220_done)
  );
  
  std_reg #(1) par_done_reg221 (
      .in(par_done_reg221_in),
      .write_en(par_done_reg221_write_en),
      .clk(clk),
      .out(par_done_reg221_out),
      .done(par_done_reg221_done)
  );
  
  std_reg #(1) par_done_reg222 (
      .in(par_done_reg222_in),
      .write_en(par_done_reg222_write_en),
      .clk(clk),
      .out(par_done_reg222_out),
      .done(par_done_reg222_done)
  );
  
  std_reg #(1) par_done_reg223 (
      .in(par_done_reg223_in),
      .write_en(par_done_reg223_write_en),
      .clk(clk),
      .out(par_done_reg223_out),
      .done(par_done_reg223_done)
  );
  
  std_reg #(1) par_done_reg224 (
      .in(par_done_reg224_in),
      .write_en(par_done_reg224_write_en),
      .clk(clk),
      .out(par_done_reg224_out),
      .done(par_done_reg224_done)
  );
  
  std_reg #(1) par_done_reg225 (
      .in(par_done_reg225_in),
      .write_en(par_done_reg225_write_en),
      .clk(clk),
      .out(par_done_reg225_out),
      .done(par_done_reg225_done)
  );
  
  std_reg #(1) par_done_reg226 (
      .in(par_done_reg226_in),
      .write_en(par_done_reg226_write_en),
      .clk(clk),
      .out(par_done_reg226_out),
      .done(par_done_reg226_done)
  );
  
  std_reg #(1) par_done_reg227 (
      .in(par_done_reg227_in),
      .write_en(par_done_reg227_write_en),
      .clk(clk),
      .out(par_done_reg227_out),
      .done(par_done_reg227_done)
  );
  
  std_reg #(1) par_done_reg228 (
      .in(par_done_reg228_in),
      .write_en(par_done_reg228_write_en),
      .clk(clk),
      .out(par_done_reg228_out),
      .done(par_done_reg228_done)
  );
  
  std_reg #(1) par_done_reg229 (
      .in(par_done_reg229_in),
      .write_en(par_done_reg229_write_en),
      .clk(clk),
      .out(par_done_reg229_out),
      .done(par_done_reg229_done)
  );
  
  std_reg #(1) par_done_reg230 (
      .in(par_done_reg230_in),
      .write_en(par_done_reg230_write_en),
      .clk(clk),
      .out(par_done_reg230_out),
      .done(par_done_reg230_done)
  );
  
  std_reg #(1) par_done_reg231 (
      .in(par_done_reg231_in),
      .write_en(par_done_reg231_write_en),
      .clk(clk),
      .out(par_done_reg231_out),
      .done(par_done_reg231_done)
  );
  
  std_reg #(1) par_reset14 (
      .in(par_reset14_in),
      .write_en(par_reset14_write_en),
      .clk(clk),
      .out(par_reset14_out),
      .done(par_reset14_done)
  );
  
  std_reg #(1) par_done_reg232 (
      .in(par_done_reg232_in),
      .write_en(par_done_reg232_write_en),
      .clk(clk),
      .out(par_done_reg232_out),
      .done(par_done_reg232_done)
  );
  
  std_reg #(1) par_done_reg233 (
      .in(par_done_reg233_in),
      .write_en(par_done_reg233_write_en),
      .clk(clk),
      .out(par_done_reg233_out),
      .done(par_done_reg233_done)
  );
  
  std_reg #(1) par_done_reg234 (
      .in(par_done_reg234_in),
      .write_en(par_done_reg234_write_en),
      .clk(clk),
      .out(par_done_reg234_out),
      .done(par_done_reg234_done)
  );
  
  std_reg #(1) par_done_reg235 (
      .in(par_done_reg235_in),
      .write_en(par_done_reg235_write_en),
      .clk(clk),
      .out(par_done_reg235_out),
      .done(par_done_reg235_done)
  );
  
  std_reg #(1) par_done_reg236 (
      .in(par_done_reg236_in),
      .write_en(par_done_reg236_write_en),
      .clk(clk),
      .out(par_done_reg236_out),
      .done(par_done_reg236_done)
  );
  
  std_reg #(1) par_done_reg237 (
      .in(par_done_reg237_in),
      .write_en(par_done_reg237_write_en),
      .clk(clk),
      .out(par_done_reg237_out),
      .done(par_done_reg237_done)
  );
  
  std_reg #(1) par_done_reg238 (
      .in(par_done_reg238_in),
      .write_en(par_done_reg238_write_en),
      .clk(clk),
      .out(par_done_reg238_out),
      .done(par_done_reg238_done)
  );
  
  std_reg #(1) par_done_reg239 (
      .in(par_done_reg239_in),
      .write_en(par_done_reg239_write_en),
      .clk(clk),
      .out(par_done_reg239_out),
      .done(par_done_reg239_done)
  );
  
  std_reg #(1) par_done_reg240 (
      .in(par_done_reg240_in),
      .write_en(par_done_reg240_write_en),
      .clk(clk),
      .out(par_done_reg240_out),
      .done(par_done_reg240_done)
  );
  
  std_reg #(1) par_done_reg241 (
      .in(par_done_reg241_in),
      .write_en(par_done_reg241_write_en),
      .clk(clk),
      .out(par_done_reg241_out),
      .done(par_done_reg241_done)
  );
  
  std_reg #(1) par_done_reg242 (
      .in(par_done_reg242_in),
      .write_en(par_done_reg242_write_en),
      .clk(clk),
      .out(par_done_reg242_out),
      .done(par_done_reg242_done)
  );
  
  std_reg #(1) par_done_reg243 (
      .in(par_done_reg243_in),
      .write_en(par_done_reg243_write_en),
      .clk(clk),
      .out(par_done_reg243_out),
      .done(par_done_reg243_done)
  );
  
  std_reg #(1) par_done_reg244 (
      .in(par_done_reg244_in),
      .write_en(par_done_reg244_write_en),
      .clk(clk),
      .out(par_done_reg244_out),
      .done(par_done_reg244_done)
  );
  
  std_reg #(1) par_done_reg245 (
      .in(par_done_reg245_in),
      .write_en(par_done_reg245_write_en),
      .clk(clk),
      .out(par_done_reg245_out),
      .done(par_done_reg245_done)
  );
  
  std_reg #(1) par_done_reg246 (
      .in(par_done_reg246_in),
      .write_en(par_done_reg246_write_en),
      .clk(clk),
      .out(par_done_reg246_out),
      .done(par_done_reg246_done)
  );
  
  std_reg #(1) par_done_reg247 (
      .in(par_done_reg247_in),
      .write_en(par_done_reg247_write_en),
      .clk(clk),
      .out(par_done_reg247_out),
      .done(par_done_reg247_done)
  );
  
  std_reg #(1) par_done_reg248 (
      .in(par_done_reg248_in),
      .write_en(par_done_reg248_write_en),
      .clk(clk),
      .out(par_done_reg248_out),
      .done(par_done_reg248_done)
  );
  
  std_reg #(1) par_done_reg249 (
      .in(par_done_reg249_in),
      .write_en(par_done_reg249_write_en),
      .clk(clk),
      .out(par_done_reg249_out),
      .done(par_done_reg249_done)
  );
  
  std_reg #(1) par_done_reg250 (
      .in(par_done_reg250_in),
      .write_en(par_done_reg250_write_en),
      .clk(clk),
      .out(par_done_reg250_out),
      .done(par_done_reg250_done)
  );
  
  std_reg #(1) par_done_reg251 (
      .in(par_done_reg251_in),
      .write_en(par_done_reg251_write_en),
      .clk(clk),
      .out(par_done_reg251_out),
      .done(par_done_reg251_done)
  );
  
  std_reg #(1) par_done_reg252 (
      .in(par_done_reg252_in),
      .write_en(par_done_reg252_write_en),
      .clk(clk),
      .out(par_done_reg252_out),
      .done(par_done_reg252_done)
  );
  
  std_reg #(1) par_done_reg253 (
      .in(par_done_reg253_in),
      .write_en(par_done_reg253_write_en),
      .clk(clk),
      .out(par_done_reg253_out),
      .done(par_done_reg253_done)
  );
  
  std_reg #(1) par_done_reg254 (
      .in(par_done_reg254_in),
      .write_en(par_done_reg254_write_en),
      .clk(clk),
      .out(par_done_reg254_out),
      .done(par_done_reg254_done)
  );
  
  std_reg #(1) par_done_reg255 (
      .in(par_done_reg255_in),
      .write_en(par_done_reg255_write_en),
      .clk(clk),
      .out(par_done_reg255_out),
      .done(par_done_reg255_done)
  );
  
  std_reg #(1) par_done_reg256 (
      .in(par_done_reg256_in),
      .write_en(par_done_reg256_write_en),
      .clk(clk),
      .out(par_done_reg256_out),
      .done(par_done_reg256_done)
  );
  
  std_reg #(1) par_done_reg257 (
      .in(par_done_reg257_in),
      .write_en(par_done_reg257_write_en),
      .clk(clk),
      .out(par_done_reg257_out),
      .done(par_done_reg257_done)
  );
  
  std_reg #(1) par_done_reg258 (
      .in(par_done_reg258_in),
      .write_en(par_done_reg258_write_en),
      .clk(clk),
      .out(par_done_reg258_out),
      .done(par_done_reg258_done)
  );
  
  std_reg #(1) par_done_reg259 (
      .in(par_done_reg259_in),
      .write_en(par_done_reg259_write_en),
      .clk(clk),
      .out(par_done_reg259_out),
      .done(par_done_reg259_done)
  );
  
  std_reg #(1) par_done_reg260 (
      .in(par_done_reg260_in),
      .write_en(par_done_reg260_write_en),
      .clk(clk),
      .out(par_done_reg260_out),
      .done(par_done_reg260_done)
  );
  
  std_reg #(1) par_done_reg261 (
      .in(par_done_reg261_in),
      .write_en(par_done_reg261_write_en),
      .clk(clk),
      .out(par_done_reg261_out),
      .done(par_done_reg261_done)
  );
  
  std_reg #(1) par_done_reg262 (
      .in(par_done_reg262_in),
      .write_en(par_done_reg262_write_en),
      .clk(clk),
      .out(par_done_reg262_out),
      .done(par_done_reg262_done)
  );
  
  std_reg #(1) par_done_reg263 (
      .in(par_done_reg263_in),
      .write_en(par_done_reg263_write_en),
      .clk(clk),
      .out(par_done_reg263_out),
      .done(par_done_reg263_done)
  );
  
  std_reg #(1) par_done_reg264 (
      .in(par_done_reg264_in),
      .write_en(par_done_reg264_write_en),
      .clk(clk),
      .out(par_done_reg264_out),
      .done(par_done_reg264_done)
  );
  
  std_reg #(1) par_done_reg265 (
      .in(par_done_reg265_in),
      .write_en(par_done_reg265_write_en),
      .clk(clk),
      .out(par_done_reg265_out),
      .done(par_done_reg265_done)
  );
  
  std_reg #(1) par_done_reg266 (
      .in(par_done_reg266_in),
      .write_en(par_done_reg266_write_en),
      .clk(clk),
      .out(par_done_reg266_out),
      .done(par_done_reg266_done)
  );
  
  std_reg #(1) par_done_reg267 (
      .in(par_done_reg267_in),
      .write_en(par_done_reg267_write_en),
      .clk(clk),
      .out(par_done_reg267_out),
      .done(par_done_reg267_done)
  );
  
  std_reg #(1) par_done_reg268 (
      .in(par_done_reg268_in),
      .write_en(par_done_reg268_write_en),
      .clk(clk),
      .out(par_done_reg268_out),
      .done(par_done_reg268_done)
  );
  
  std_reg #(1) par_done_reg269 (
      .in(par_done_reg269_in),
      .write_en(par_done_reg269_write_en),
      .clk(clk),
      .out(par_done_reg269_out),
      .done(par_done_reg269_done)
  );
  
  std_reg #(1) par_done_reg270 (
      .in(par_done_reg270_in),
      .write_en(par_done_reg270_write_en),
      .clk(clk),
      .out(par_done_reg270_out),
      .done(par_done_reg270_done)
  );
  
  std_reg #(1) par_done_reg271 (
      .in(par_done_reg271_in),
      .write_en(par_done_reg271_write_en),
      .clk(clk),
      .out(par_done_reg271_out),
      .done(par_done_reg271_done)
  );
  
  std_reg #(1) par_done_reg272 (
      .in(par_done_reg272_in),
      .write_en(par_done_reg272_write_en),
      .clk(clk),
      .out(par_done_reg272_out),
      .done(par_done_reg272_done)
  );
  
  std_reg #(1) par_done_reg273 (
      .in(par_done_reg273_in),
      .write_en(par_done_reg273_write_en),
      .clk(clk),
      .out(par_done_reg273_out),
      .done(par_done_reg273_done)
  );
  
  std_reg #(1) par_done_reg274 (
      .in(par_done_reg274_in),
      .write_en(par_done_reg274_write_en),
      .clk(clk),
      .out(par_done_reg274_out),
      .done(par_done_reg274_done)
  );
  
  std_reg #(1) par_done_reg275 (
      .in(par_done_reg275_in),
      .write_en(par_done_reg275_write_en),
      .clk(clk),
      .out(par_done_reg275_out),
      .done(par_done_reg275_done)
  );
  
  std_reg #(1) par_done_reg276 (
      .in(par_done_reg276_in),
      .write_en(par_done_reg276_write_en),
      .clk(clk),
      .out(par_done_reg276_out),
      .done(par_done_reg276_done)
  );
  
  std_reg #(1) par_done_reg277 (
      .in(par_done_reg277_in),
      .write_en(par_done_reg277_write_en),
      .clk(clk),
      .out(par_done_reg277_out),
      .done(par_done_reg277_done)
  );
  
  std_reg #(1) par_done_reg278 (
      .in(par_done_reg278_in),
      .write_en(par_done_reg278_write_en),
      .clk(clk),
      .out(par_done_reg278_out),
      .done(par_done_reg278_done)
  );
  
  std_reg #(1) par_done_reg279 (
      .in(par_done_reg279_in),
      .write_en(par_done_reg279_write_en),
      .clk(clk),
      .out(par_done_reg279_out),
      .done(par_done_reg279_done)
  );
  
  std_reg #(1) par_done_reg280 (
      .in(par_done_reg280_in),
      .write_en(par_done_reg280_write_en),
      .clk(clk),
      .out(par_done_reg280_out),
      .done(par_done_reg280_done)
  );
  
  std_reg #(1) par_done_reg281 (
      .in(par_done_reg281_in),
      .write_en(par_done_reg281_write_en),
      .clk(clk),
      .out(par_done_reg281_out),
      .done(par_done_reg281_done)
  );
  
  std_reg #(1) par_reset15 (
      .in(par_reset15_in),
      .write_en(par_reset15_write_en),
      .clk(clk),
      .out(par_reset15_out),
      .done(par_reset15_done)
  );
  
  std_reg #(1) par_done_reg282 (
      .in(par_done_reg282_in),
      .write_en(par_done_reg282_write_en),
      .clk(clk),
      .out(par_done_reg282_out),
      .done(par_done_reg282_done)
  );
  
  std_reg #(1) par_done_reg283 (
      .in(par_done_reg283_in),
      .write_en(par_done_reg283_write_en),
      .clk(clk),
      .out(par_done_reg283_out),
      .done(par_done_reg283_done)
  );
  
  std_reg #(1) par_done_reg284 (
      .in(par_done_reg284_in),
      .write_en(par_done_reg284_write_en),
      .clk(clk),
      .out(par_done_reg284_out),
      .done(par_done_reg284_done)
  );
  
  std_reg #(1) par_done_reg285 (
      .in(par_done_reg285_in),
      .write_en(par_done_reg285_write_en),
      .clk(clk),
      .out(par_done_reg285_out),
      .done(par_done_reg285_done)
  );
  
  std_reg #(1) par_done_reg286 (
      .in(par_done_reg286_in),
      .write_en(par_done_reg286_write_en),
      .clk(clk),
      .out(par_done_reg286_out),
      .done(par_done_reg286_done)
  );
  
  std_reg #(1) par_done_reg287 (
      .in(par_done_reg287_in),
      .write_en(par_done_reg287_write_en),
      .clk(clk),
      .out(par_done_reg287_out),
      .done(par_done_reg287_done)
  );
  
  std_reg #(1) par_done_reg288 (
      .in(par_done_reg288_in),
      .write_en(par_done_reg288_write_en),
      .clk(clk),
      .out(par_done_reg288_out),
      .done(par_done_reg288_done)
  );
  
  std_reg #(1) par_done_reg289 (
      .in(par_done_reg289_in),
      .write_en(par_done_reg289_write_en),
      .clk(clk),
      .out(par_done_reg289_out),
      .done(par_done_reg289_done)
  );
  
  std_reg #(1) par_done_reg290 (
      .in(par_done_reg290_in),
      .write_en(par_done_reg290_write_en),
      .clk(clk),
      .out(par_done_reg290_out),
      .done(par_done_reg290_done)
  );
  
  std_reg #(1) par_done_reg291 (
      .in(par_done_reg291_in),
      .write_en(par_done_reg291_write_en),
      .clk(clk),
      .out(par_done_reg291_out),
      .done(par_done_reg291_done)
  );
  
  std_reg #(1) par_done_reg292 (
      .in(par_done_reg292_in),
      .write_en(par_done_reg292_write_en),
      .clk(clk),
      .out(par_done_reg292_out),
      .done(par_done_reg292_done)
  );
  
  std_reg #(1) par_done_reg293 (
      .in(par_done_reg293_in),
      .write_en(par_done_reg293_write_en),
      .clk(clk),
      .out(par_done_reg293_out),
      .done(par_done_reg293_done)
  );
  
  std_reg #(1) par_done_reg294 (
      .in(par_done_reg294_in),
      .write_en(par_done_reg294_write_en),
      .clk(clk),
      .out(par_done_reg294_out),
      .done(par_done_reg294_done)
  );
  
  std_reg #(1) par_done_reg295 (
      .in(par_done_reg295_in),
      .write_en(par_done_reg295_write_en),
      .clk(clk),
      .out(par_done_reg295_out),
      .done(par_done_reg295_done)
  );
  
  std_reg #(1) par_done_reg296 (
      .in(par_done_reg296_in),
      .write_en(par_done_reg296_write_en),
      .clk(clk),
      .out(par_done_reg296_out),
      .done(par_done_reg296_done)
  );
  
  std_reg #(1) par_done_reg297 (
      .in(par_done_reg297_in),
      .write_en(par_done_reg297_write_en),
      .clk(clk),
      .out(par_done_reg297_out),
      .done(par_done_reg297_done)
  );
  
  std_reg #(1) par_done_reg298 (
      .in(par_done_reg298_in),
      .write_en(par_done_reg298_write_en),
      .clk(clk),
      .out(par_done_reg298_out),
      .done(par_done_reg298_done)
  );
  
  std_reg #(1) par_done_reg299 (
      .in(par_done_reg299_in),
      .write_en(par_done_reg299_write_en),
      .clk(clk),
      .out(par_done_reg299_out),
      .done(par_done_reg299_done)
  );
  
  std_reg #(1) par_done_reg300 (
      .in(par_done_reg300_in),
      .write_en(par_done_reg300_write_en),
      .clk(clk),
      .out(par_done_reg300_out),
      .done(par_done_reg300_done)
  );
  
  std_reg #(1) par_done_reg301 (
      .in(par_done_reg301_in),
      .write_en(par_done_reg301_write_en),
      .clk(clk),
      .out(par_done_reg301_out),
      .done(par_done_reg301_done)
  );
  
  std_reg #(1) par_done_reg302 (
      .in(par_done_reg302_in),
      .write_en(par_done_reg302_write_en),
      .clk(clk),
      .out(par_done_reg302_out),
      .done(par_done_reg302_done)
  );
  
  std_reg #(1) par_done_reg303 (
      .in(par_done_reg303_in),
      .write_en(par_done_reg303_write_en),
      .clk(clk),
      .out(par_done_reg303_out),
      .done(par_done_reg303_done)
  );
  
  std_reg #(1) par_done_reg304 (
      .in(par_done_reg304_in),
      .write_en(par_done_reg304_write_en),
      .clk(clk),
      .out(par_done_reg304_out),
      .done(par_done_reg304_done)
  );
  
  std_reg #(1) par_done_reg305 (
      .in(par_done_reg305_in),
      .write_en(par_done_reg305_write_en),
      .clk(clk),
      .out(par_done_reg305_out),
      .done(par_done_reg305_done)
  );
  
  std_reg #(1) par_done_reg306 (
      .in(par_done_reg306_in),
      .write_en(par_done_reg306_write_en),
      .clk(clk),
      .out(par_done_reg306_out),
      .done(par_done_reg306_done)
  );
  
  std_reg #(1) par_done_reg307 (
      .in(par_done_reg307_in),
      .write_en(par_done_reg307_write_en),
      .clk(clk),
      .out(par_done_reg307_out),
      .done(par_done_reg307_done)
  );
  
  std_reg #(1) par_done_reg308 (
      .in(par_done_reg308_in),
      .write_en(par_done_reg308_write_en),
      .clk(clk),
      .out(par_done_reg308_out),
      .done(par_done_reg308_done)
  );
  
  std_reg #(1) par_done_reg309 (
      .in(par_done_reg309_in),
      .write_en(par_done_reg309_write_en),
      .clk(clk),
      .out(par_done_reg309_out),
      .done(par_done_reg309_done)
  );
  
  std_reg #(1) par_done_reg310 (
      .in(par_done_reg310_in),
      .write_en(par_done_reg310_write_en),
      .clk(clk),
      .out(par_done_reg310_out),
      .done(par_done_reg310_done)
  );
  
  std_reg #(1) par_done_reg311 (
      .in(par_done_reg311_in),
      .write_en(par_done_reg311_write_en),
      .clk(clk),
      .out(par_done_reg311_out),
      .done(par_done_reg311_done)
  );
  
  std_reg #(1) par_done_reg312 (
      .in(par_done_reg312_in),
      .write_en(par_done_reg312_write_en),
      .clk(clk),
      .out(par_done_reg312_out),
      .done(par_done_reg312_done)
  );
  
  std_reg #(1) par_done_reg313 (
      .in(par_done_reg313_in),
      .write_en(par_done_reg313_write_en),
      .clk(clk),
      .out(par_done_reg313_out),
      .done(par_done_reg313_done)
  );
  
  std_reg #(1) par_done_reg314 (
      .in(par_done_reg314_in),
      .write_en(par_done_reg314_write_en),
      .clk(clk),
      .out(par_done_reg314_out),
      .done(par_done_reg314_done)
  );
  
  std_reg #(1) par_reset16 (
      .in(par_reset16_in),
      .write_en(par_reset16_write_en),
      .clk(clk),
      .out(par_reset16_out),
      .done(par_reset16_done)
  );
  
  std_reg #(1) par_done_reg315 (
      .in(par_done_reg315_in),
      .write_en(par_done_reg315_write_en),
      .clk(clk),
      .out(par_done_reg315_out),
      .done(par_done_reg315_done)
  );
  
  std_reg #(1) par_done_reg316 (
      .in(par_done_reg316_in),
      .write_en(par_done_reg316_write_en),
      .clk(clk),
      .out(par_done_reg316_out),
      .done(par_done_reg316_done)
  );
  
  std_reg #(1) par_done_reg317 (
      .in(par_done_reg317_in),
      .write_en(par_done_reg317_write_en),
      .clk(clk),
      .out(par_done_reg317_out),
      .done(par_done_reg317_done)
  );
  
  std_reg #(1) par_done_reg318 (
      .in(par_done_reg318_in),
      .write_en(par_done_reg318_write_en),
      .clk(clk),
      .out(par_done_reg318_out),
      .done(par_done_reg318_done)
  );
  
  std_reg #(1) par_done_reg319 (
      .in(par_done_reg319_in),
      .write_en(par_done_reg319_write_en),
      .clk(clk),
      .out(par_done_reg319_out),
      .done(par_done_reg319_done)
  );
  
  std_reg #(1) par_done_reg320 (
      .in(par_done_reg320_in),
      .write_en(par_done_reg320_write_en),
      .clk(clk),
      .out(par_done_reg320_out),
      .done(par_done_reg320_done)
  );
  
  std_reg #(1) par_done_reg321 (
      .in(par_done_reg321_in),
      .write_en(par_done_reg321_write_en),
      .clk(clk),
      .out(par_done_reg321_out),
      .done(par_done_reg321_done)
  );
  
  std_reg #(1) par_done_reg322 (
      .in(par_done_reg322_in),
      .write_en(par_done_reg322_write_en),
      .clk(clk),
      .out(par_done_reg322_out),
      .done(par_done_reg322_done)
  );
  
  std_reg #(1) par_done_reg323 (
      .in(par_done_reg323_in),
      .write_en(par_done_reg323_write_en),
      .clk(clk),
      .out(par_done_reg323_out),
      .done(par_done_reg323_done)
  );
  
  std_reg #(1) par_done_reg324 (
      .in(par_done_reg324_in),
      .write_en(par_done_reg324_write_en),
      .clk(clk),
      .out(par_done_reg324_out),
      .done(par_done_reg324_done)
  );
  
  std_reg #(1) par_done_reg325 (
      .in(par_done_reg325_in),
      .write_en(par_done_reg325_write_en),
      .clk(clk),
      .out(par_done_reg325_out),
      .done(par_done_reg325_done)
  );
  
  std_reg #(1) par_done_reg326 (
      .in(par_done_reg326_in),
      .write_en(par_done_reg326_write_en),
      .clk(clk),
      .out(par_done_reg326_out),
      .done(par_done_reg326_done)
  );
  
  std_reg #(1) par_done_reg327 (
      .in(par_done_reg327_in),
      .write_en(par_done_reg327_write_en),
      .clk(clk),
      .out(par_done_reg327_out),
      .done(par_done_reg327_done)
  );
  
  std_reg #(1) par_done_reg328 (
      .in(par_done_reg328_in),
      .write_en(par_done_reg328_write_en),
      .clk(clk),
      .out(par_done_reg328_out),
      .done(par_done_reg328_done)
  );
  
  std_reg #(1) par_done_reg329 (
      .in(par_done_reg329_in),
      .write_en(par_done_reg329_write_en),
      .clk(clk),
      .out(par_done_reg329_out),
      .done(par_done_reg329_done)
  );
  
  std_reg #(1) par_done_reg330 (
      .in(par_done_reg330_in),
      .write_en(par_done_reg330_write_en),
      .clk(clk),
      .out(par_done_reg330_out),
      .done(par_done_reg330_done)
  );
  
  std_reg #(1) par_done_reg331 (
      .in(par_done_reg331_in),
      .write_en(par_done_reg331_write_en),
      .clk(clk),
      .out(par_done_reg331_out),
      .done(par_done_reg331_done)
  );
  
  std_reg #(1) par_done_reg332 (
      .in(par_done_reg332_in),
      .write_en(par_done_reg332_write_en),
      .clk(clk),
      .out(par_done_reg332_out),
      .done(par_done_reg332_done)
  );
  
  std_reg #(1) par_done_reg333 (
      .in(par_done_reg333_in),
      .write_en(par_done_reg333_write_en),
      .clk(clk),
      .out(par_done_reg333_out),
      .done(par_done_reg333_done)
  );
  
  std_reg #(1) par_done_reg334 (
      .in(par_done_reg334_in),
      .write_en(par_done_reg334_write_en),
      .clk(clk),
      .out(par_done_reg334_out),
      .done(par_done_reg334_done)
  );
  
  std_reg #(1) par_done_reg335 (
      .in(par_done_reg335_in),
      .write_en(par_done_reg335_write_en),
      .clk(clk),
      .out(par_done_reg335_out),
      .done(par_done_reg335_done)
  );
  
  std_reg #(1) par_done_reg336 (
      .in(par_done_reg336_in),
      .write_en(par_done_reg336_write_en),
      .clk(clk),
      .out(par_done_reg336_out),
      .done(par_done_reg336_done)
  );
  
  std_reg #(1) par_done_reg337 (
      .in(par_done_reg337_in),
      .write_en(par_done_reg337_write_en),
      .clk(clk),
      .out(par_done_reg337_out),
      .done(par_done_reg337_done)
  );
  
  std_reg #(1) par_done_reg338 (
      .in(par_done_reg338_in),
      .write_en(par_done_reg338_write_en),
      .clk(clk),
      .out(par_done_reg338_out),
      .done(par_done_reg338_done)
  );
  
  std_reg #(1) par_done_reg339 (
      .in(par_done_reg339_in),
      .write_en(par_done_reg339_write_en),
      .clk(clk),
      .out(par_done_reg339_out),
      .done(par_done_reg339_done)
  );
  
  std_reg #(1) par_done_reg340 (
      .in(par_done_reg340_in),
      .write_en(par_done_reg340_write_en),
      .clk(clk),
      .out(par_done_reg340_out),
      .done(par_done_reg340_done)
  );
  
  std_reg #(1) par_done_reg341 (
      .in(par_done_reg341_in),
      .write_en(par_done_reg341_write_en),
      .clk(clk),
      .out(par_done_reg341_out),
      .done(par_done_reg341_done)
  );
  
  std_reg #(1) par_done_reg342 (
      .in(par_done_reg342_in),
      .write_en(par_done_reg342_write_en),
      .clk(clk),
      .out(par_done_reg342_out),
      .done(par_done_reg342_done)
  );
  
  std_reg #(1) par_done_reg343 (
      .in(par_done_reg343_in),
      .write_en(par_done_reg343_write_en),
      .clk(clk),
      .out(par_done_reg343_out),
      .done(par_done_reg343_done)
  );
  
  std_reg #(1) par_done_reg344 (
      .in(par_done_reg344_in),
      .write_en(par_done_reg344_write_en),
      .clk(clk),
      .out(par_done_reg344_out),
      .done(par_done_reg344_done)
  );
  
  std_reg #(1) par_done_reg345 (
      .in(par_done_reg345_in),
      .write_en(par_done_reg345_write_en),
      .clk(clk),
      .out(par_done_reg345_out),
      .done(par_done_reg345_done)
  );
  
  std_reg #(1) par_done_reg346 (
      .in(par_done_reg346_in),
      .write_en(par_done_reg346_write_en),
      .clk(clk),
      .out(par_done_reg346_out),
      .done(par_done_reg346_done)
  );
  
  std_reg #(1) par_done_reg347 (
      .in(par_done_reg347_in),
      .write_en(par_done_reg347_write_en),
      .clk(clk),
      .out(par_done_reg347_out),
      .done(par_done_reg347_done)
  );
  
  std_reg #(1) par_done_reg348 (
      .in(par_done_reg348_in),
      .write_en(par_done_reg348_write_en),
      .clk(clk),
      .out(par_done_reg348_out),
      .done(par_done_reg348_done)
  );
  
  std_reg #(1) par_done_reg349 (
      .in(par_done_reg349_in),
      .write_en(par_done_reg349_write_en),
      .clk(clk),
      .out(par_done_reg349_out),
      .done(par_done_reg349_done)
  );
  
  std_reg #(1) par_done_reg350 (
      .in(par_done_reg350_in),
      .write_en(par_done_reg350_write_en),
      .clk(clk),
      .out(par_done_reg350_out),
      .done(par_done_reg350_done)
  );
  
  std_reg #(1) par_done_reg351 (
      .in(par_done_reg351_in),
      .write_en(par_done_reg351_write_en),
      .clk(clk),
      .out(par_done_reg351_out),
      .done(par_done_reg351_done)
  );
  
  std_reg #(1) par_done_reg352 (
      .in(par_done_reg352_in),
      .write_en(par_done_reg352_write_en),
      .clk(clk),
      .out(par_done_reg352_out),
      .done(par_done_reg352_done)
  );
  
  std_reg #(1) par_done_reg353 (
      .in(par_done_reg353_in),
      .write_en(par_done_reg353_write_en),
      .clk(clk),
      .out(par_done_reg353_out),
      .done(par_done_reg353_done)
  );
  
  std_reg #(1) par_done_reg354 (
      .in(par_done_reg354_in),
      .write_en(par_done_reg354_write_en),
      .clk(clk),
      .out(par_done_reg354_out),
      .done(par_done_reg354_done)
  );
  
  std_reg #(1) par_done_reg355 (
      .in(par_done_reg355_in),
      .write_en(par_done_reg355_write_en),
      .clk(clk),
      .out(par_done_reg355_out),
      .done(par_done_reg355_done)
  );
  
  std_reg #(1) par_done_reg356 (
      .in(par_done_reg356_in),
      .write_en(par_done_reg356_write_en),
      .clk(clk),
      .out(par_done_reg356_out),
      .done(par_done_reg356_done)
  );
  
  std_reg #(1) par_done_reg357 (
      .in(par_done_reg357_in),
      .write_en(par_done_reg357_write_en),
      .clk(clk),
      .out(par_done_reg357_out),
      .done(par_done_reg357_done)
  );
  
  std_reg #(1) par_done_reg358 (
      .in(par_done_reg358_in),
      .write_en(par_done_reg358_write_en),
      .clk(clk),
      .out(par_done_reg358_out),
      .done(par_done_reg358_done)
  );
  
  std_reg #(1) par_done_reg359 (
      .in(par_done_reg359_in),
      .write_en(par_done_reg359_write_en),
      .clk(clk),
      .out(par_done_reg359_out),
      .done(par_done_reg359_done)
  );
  
  std_reg #(1) par_done_reg360 (
      .in(par_done_reg360_in),
      .write_en(par_done_reg360_write_en),
      .clk(clk),
      .out(par_done_reg360_out),
      .done(par_done_reg360_done)
  );
  
  std_reg #(1) par_done_reg361 (
      .in(par_done_reg361_in),
      .write_en(par_done_reg361_write_en),
      .clk(clk),
      .out(par_done_reg361_out),
      .done(par_done_reg361_done)
  );
  
  std_reg #(1) par_done_reg362 (
      .in(par_done_reg362_in),
      .write_en(par_done_reg362_write_en),
      .clk(clk),
      .out(par_done_reg362_out),
      .done(par_done_reg362_done)
  );
  
  std_reg #(1) par_done_reg363 (
      .in(par_done_reg363_in),
      .write_en(par_done_reg363_write_en),
      .clk(clk),
      .out(par_done_reg363_out),
      .done(par_done_reg363_done)
  );
  
  std_reg #(1) par_done_reg364 (
      .in(par_done_reg364_in),
      .write_en(par_done_reg364_write_en),
      .clk(clk),
      .out(par_done_reg364_out),
      .done(par_done_reg364_done)
  );
  
  std_reg #(1) par_done_reg365 (
      .in(par_done_reg365_in),
      .write_en(par_done_reg365_write_en),
      .clk(clk),
      .out(par_done_reg365_out),
      .done(par_done_reg365_done)
  );
  
  std_reg #(1) par_done_reg366 (
      .in(par_done_reg366_in),
      .write_en(par_done_reg366_write_en),
      .clk(clk),
      .out(par_done_reg366_out),
      .done(par_done_reg366_done)
  );
  
  std_reg #(1) par_done_reg367 (
      .in(par_done_reg367_in),
      .write_en(par_done_reg367_write_en),
      .clk(clk),
      .out(par_done_reg367_out),
      .done(par_done_reg367_done)
  );
  
  std_reg #(1) par_done_reg368 (
      .in(par_done_reg368_in),
      .write_en(par_done_reg368_write_en),
      .clk(clk),
      .out(par_done_reg368_out),
      .done(par_done_reg368_done)
  );
  
  std_reg #(1) par_reset17 (
      .in(par_reset17_in),
      .write_en(par_reset17_write_en),
      .clk(clk),
      .out(par_reset17_out),
      .done(par_reset17_done)
  );
  
  std_reg #(1) par_done_reg369 (
      .in(par_done_reg369_in),
      .write_en(par_done_reg369_write_en),
      .clk(clk),
      .out(par_done_reg369_out),
      .done(par_done_reg369_done)
  );
  
  std_reg #(1) par_done_reg370 (
      .in(par_done_reg370_in),
      .write_en(par_done_reg370_write_en),
      .clk(clk),
      .out(par_done_reg370_out),
      .done(par_done_reg370_done)
  );
  
  std_reg #(1) par_done_reg371 (
      .in(par_done_reg371_in),
      .write_en(par_done_reg371_write_en),
      .clk(clk),
      .out(par_done_reg371_out),
      .done(par_done_reg371_done)
  );
  
  std_reg #(1) par_done_reg372 (
      .in(par_done_reg372_in),
      .write_en(par_done_reg372_write_en),
      .clk(clk),
      .out(par_done_reg372_out),
      .done(par_done_reg372_done)
  );
  
  std_reg #(1) par_done_reg373 (
      .in(par_done_reg373_in),
      .write_en(par_done_reg373_write_en),
      .clk(clk),
      .out(par_done_reg373_out),
      .done(par_done_reg373_done)
  );
  
  std_reg #(1) par_done_reg374 (
      .in(par_done_reg374_in),
      .write_en(par_done_reg374_write_en),
      .clk(clk),
      .out(par_done_reg374_out),
      .done(par_done_reg374_done)
  );
  
  std_reg #(1) par_done_reg375 (
      .in(par_done_reg375_in),
      .write_en(par_done_reg375_write_en),
      .clk(clk),
      .out(par_done_reg375_out),
      .done(par_done_reg375_done)
  );
  
  std_reg #(1) par_done_reg376 (
      .in(par_done_reg376_in),
      .write_en(par_done_reg376_write_en),
      .clk(clk),
      .out(par_done_reg376_out),
      .done(par_done_reg376_done)
  );
  
  std_reg #(1) par_done_reg377 (
      .in(par_done_reg377_in),
      .write_en(par_done_reg377_write_en),
      .clk(clk),
      .out(par_done_reg377_out),
      .done(par_done_reg377_done)
  );
  
  std_reg #(1) par_done_reg378 (
      .in(par_done_reg378_in),
      .write_en(par_done_reg378_write_en),
      .clk(clk),
      .out(par_done_reg378_out),
      .done(par_done_reg378_done)
  );
  
  std_reg #(1) par_done_reg379 (
      .in(par_done_reg379_in),
      .write_en(par_done_reg379_write_en),
      .clk(clk),
      .out(par_done_reg379_out),
      .done(par_done_reg379_done)
  );
  
  std_reg #(1) par_done_reg380 (
      .in(par_done_reg380_in),
      .write_en(par_done_reg380_write_en),
      .clk(clk),
      .out(par_done_reg380_out),
      .done(par_done_reg380_done)
  );
  
  std_reg #(1) par_done_reg381 (
      .in(par_done_reg381_in),
      .write_en(par_done_reg381_write_en),
      .clk(clk),
      .out(par_done_reg381_out),
      .done(par_done_reg381_done)
  );
  
  std_reg #(1) par_done_reg382 (
      .in(par_done_reg382_in),
      .write_en(par_done_reg382_write_en),
      .clk(clk),
      .out(par_done_reg382_out),
      .done(par_done_reg382_done)
  );
  
  std_reg #(1) par_done_reg383 (
      .in(par_done_reg383_in),
      .write_en(par_done_reg383_write_en),
      .clk(clk),
      .out(par_done_reg383_out),
      .done(par_done_reg383_done)
  );
  
  std_reg #(1) par_done_reg384 (
      .in(par_done_reg384_in),
      .write_en(par_done_reg384_write_en),
      .clk(clk),
      .out(par_done_reg384_out),
      .done(par_done_reg384_done)
  );
  
  std_reg #(1) par_done_reg385 (
      .in(par_done_reg385_in),
      .write_en(par_done_reg385_write_en),
      .clk(clk),
      .out(par_done_reg385_out),
      .done(par_done_reg385_done)
  );
  
  std_reg #(1) par_done_reg386 (
      .in(par_done_reg386_in),
      .write_en(par_done_reg386_write_en),
      .clk(clk),
      .out(par_done_reg386_out),
      .done(par_done_reg386_done)
  );
  
  std_reg #(1) par_done_reg387 (
      .in(par_done_reg387_in),
      .write_en(par_done_reg387_write_en),
      .clk(clk),
      .out(par_done_reg387_out),
      .done(par_done_reg387_done)
  );
  
  std_reg #(1) par_done_reg388 (
      .in(par_done_reg388_in),
      .write_en(par_done_reg388_write_en),
      .clk(clk),
      .out(par_done_reg388_out),
      .done(par_done_reg388_done)
  );
  
  std_reg #(1) par_done_reg389 (
      .in(par_done_reg389_in),
      .write_en(par_done_reg389_write_en),
      .clk(clk),
      .out(par_done_reg389_out),
      .done(par_done_reg389_done)
  );
  
  std_reg #(1) par_done_reg390 (
      .in(par_done_reg390_in),
      .write_en(par_done_reg390_write_en),
      .clk(clk),
      .out(par_done_reg390_out),
      .done(par_done_reg390_done)
  );
  
  std_reg #(1) par_done_reg391 (
      .in(par_done_reg391_in),
      .write_en(par_done_reg391_write_en),
      .clk(clk),
      .out(par_done_reg391_out),
      .done(par_done_reg391_done)
  );
  
  std_reg #(1) par_done_reg392 (
      .in(par_done_reg392_in),
      .write_en(par_done_reg392_write_en),
      .clk(clk),
      .out(par_done_reg392_out),
      .done(par_done_reg392_done)
  );
  
  std_reg #(1) par_done_reg393 (
      .in(par_done_reg393_in),
      .write_en(par_done_reg393_write_en),
      .clk(clk),
      .out(par_done_reg393_out),
      .done(par_done_reg393_done)
  );
  
  std_reg #(1) par_done_reg394 (
      .in(par_done_reg394_in),
      .write_en(par_done_reg394_write_en),
      .clk(clk),
      .out(par_done_reg394_out),
      .done(par_done_reg394_done)
  );
  
  std_reg #(1) par_done_reg395 (
      .in(par_done_reg395_in),
      .write_en(par_done_reg395_write_en),
      .clk(clk),
      .out(par_done_reg395_out),
      .done(par_done_reg395_done)
  );
  
  std_reg #(1) par_done_reg396 (
      .in(par_done_reg396_in),
      .write_en(par_done_reg396_write_en),
      .clk(clk),
      .out(par_done_reg396_out),
      .done(par_done_reg396_done)
  );
  
  std_reg #(1) par_done_reg397 (
      .in(par_done_reg397_in),
      .write_en(par_done_reg397_write_en),
      .clk(clk),
      .out(par_done_reg397_out),
      .done(par_done_reg397_done)
  );
  
  std_reg #(1) par_done_reg398 (
      .in(par_done_reg398_in),
      .write_en(par_done_reg398_write_en),
      .clk(clk),
      .out(par_done_reg398_out),
      .done(par_done_reg398_done)
  );
  
  std_reg #(1) par_done_reg399 (
      .in(par_done_reg399_in),
      .write_en(par_done_reg399_write_en),
      .clk(clk),
      .out(par_done_reg399_out),
      .done(par_done_reg399_done)
  );
  
  std_reg #(1) par_done_reg400 (
      .in(par_done_reg400_in),
      .write_en(par_done_reg400_write_en),
      .clk(clk),
      .out(par_done_reg400_out),
      .done(par_done_reg400_done)
  );
  
  std_reg #(1) par_done_reg401 (
      .in(par_done_reg401_in),
      .write_en(par_done_reg401_write_en),
      .clk(clk),
      .out(par_done_reg401_out),
      .done(par_done_reg401_done)
  );
  
  std_reg #(1) par_reset18 (
      .in(par_reset18_in),
      .write_en(par_reset18_write_en),
      .clk(clk),
      .out(par_reset18_out),
      .done(par_reset18_done)
  );
  
  std_reg #(1) par_done_reg402 (
      .in(par_done_reg402_in),
      .write_en(par_done_reg402_write_en),
      .clk(clk),
      .out(par_done_reg402_out),
      .done(par_done_reg402_done)
  );
  
  std_reg #(1) par_done_reg403 (
      .in(par_done_reg403_in),
      .write_en(par_done_reg403_write_en),
      .clk(clk),
      .out(par_done_reg403_out),
      .done(par_done_reg403_done)
  );
  
  std_reg #(1) par_done_reg404 (
      .in(par_done_reg404_in),
      .write_en(par_done_reg404_write_en),
      .clk(clk),
      .out(par_done_reg404_out),
      .done(par_done_reg404_done)
  );
  
  std_reg #(1) par_done_reg405 (
      .in(par_done_reg405_in),
      .write_en(par_done_reg405_write_en),
      .clk(clk),
      .out(par_done_reg405_out),
      .done(par_done_reg405_done)
  );
  
  std_reg #(1) par_done_reg406 (
      .in(par_done_reg406_in),
      .write_en(par_done_reg406_write_en),
      .clk(clk),
      .out(par_done_reg406_out),
      .done(par_done_reg406_done)
  );
  
  std_reg #(1) par_done_reg407 (
      .in(par_done_reg407_in),
      .write_en(par_done_reg407_write_en),
      .clk(clk),
      .out(par_done_reg407_out),
      .done(par_done_reg407_done)
  );
  
  std_reg #(1) par_done_reg408 (
      .in(par_done_reg408_in),
      .write_en(par_done_reg408_write_en),
      .clk(clk),
      .out(par_done_reg408_out),
      .done(par_done_reg408_done)
  );
  
  std_reg #(1) par_done_reg409 (
      .in(par_done_reg409_in),
      .write_en(par_done_reg409_write_en),
      .clk(clk),
      .out(par_done_reg409_out),
      .done(par_done_reg409_done)
  );
  
  std_reg #(1) par_done_reg410 (
      .in(par_done_reg410_in),
      .write_en(par_done_reg410_write_en),
      .clk(clk),
      .out(par_done_reg410_out),
      .done(par_done_reg410_done)
  );
  
  std_reg #(1) par_done_reg411 (
      .in(par_done_reg411_in),
      .write_en(par_done_reg411_write_en),
      .clk(clk),
      .out(par_done_reg411_out),
      .done(par_done_reg411_done)
  );
  
  std_reg #(1) par_done_reg412 (
      .in(par_done_reg412_in),
      .write_en(par_done_reg412_write_en),
      .clk(clk),
      .out(par_done_reg412_out),
      .done(par_done_reg412_done)
  );
  
  std_reg #(1) par_done_reg413 (
      .in(par_done_reg413_in),
      .write_en(par_done_reg413_write_en),
      .clk(clk),
      .out(par_done_reg413_out),
      .done(par_done_reg413_done)
  );
  
  std_reg #(1) par_done_reg414 (
      .in(par_done_reg414_in),
      .write_en(par_done_reg414_write_en),
      .clk(clk),
      .out(par_done_reg414_out),
      .done(par_done_reg414_done)
  );
  
  std_reg #(1) par_done_reg415 (
      .in(par_done_reg415_in),
      .write_en(par_done_reg415_write_en),
      .clk(clk),
      .out(par_done_reg415_out),
      .done(par_done_reg415_done)
  );
  
  std_reg #(1) par_done_reg416 (
      .in(par_done_reg416_in),
      .write_en(par_done_reg416_write_en),
      .clk(clk),
      .out(par_done_reg416_out),
      .done(par_done_reg416_done)
  );
  
  std_reg #(1) par_done_reg417 (
      .in(par_done_reg417_in),
      .write_en(par_done_reg417_write_en),
      .clk(clk),
      .out(par_done_reg417_out),
      .done(par_done_reg417_done)
  );
  
  std_reg #(1) par_done_reg418 (
      .in(par_done_reg418_in),
      .write_en(par_done_reg418_write_en),
      .clk(clk),
      .out(par_done_reg418_out),
      .done(par_done_reg418_done)
  );
  
  std_reg #(1) par_done_reg419 (
      .in(par_done_reg419_in),
      .write_en(par_done_reg419_write_en),
      .clk(clk),
      .out(par_done_reg419_out),
      .done(par_done_reg419_done)
  );
  
  std_reg #(1) par_done_reg420 (
      .in(par_done_reg420_in),
      .write_en(par_done_reg420_write_en),
      .clk(clk),
      .out(par_done_reg420_out),
      .done(par_done_reg420_done)
  );
  
  std_reg #(1) par_done_reg421 (
      .in(par_done_reg421_in),
      .write_en(par_done_reg421_write_en),
      .clk(clk),
      .out(par_done_reg421_out),
      .done(par_done_reg421_done)
  );
  
  std_reg #(1) par_done_reg422 (
      .in(par_done_reg422_in),
      .write_en(par_done_reg422_write_en),
      .clk(clk),
      .out(par_done_reg422_out),
      .done(par_done_reg422_done)
  );
  
  std_reg #(1) par_done_reg423 (
      .in(par_done_reg423_in),
      .write_en(par_done_reg423_write_en),
      .clk(clk),
      .out(par_done_reg423_out),
      .done(par_done_reg423_done)
  );
  
  std_reg #(1) par_done_reg424 (
      .in(par_done_reg424_in),
      .write_en(par_done_reg424_write_en),
      .clk(clk),
      .out(par_done_reg424_out),
      .done(par_done_reg424_done)
  );
  
  std_reg #(1) par_done_reg425 (
      .in(par_done_reg425_in),
      .write_en(par_done_reg425_write_en),
      .clk(clk),
      .out(par_done_reg425_out),
      .done(par_done_reg425_done)
  );
  
  std_reg #(1) par_done_reg426 (
      .in(par_done_reg426_in),
      .write_en(par_done_reg426_write_en),
      .clk(clk),
      .out(par_done_reg426_out),
      .done(par_done_reg426_done)
  );
  
  std_reg #(1) par_done_reg427 (
      .in(par_done_reg427_in),
      .write_en(par_done_reg427_write_en),
      .clk(clk),
      .out(par_done_reg427_out),
      .done(par_done_reg427_done)
  );
  
  std_reg #(1) par_done_reg428 (
      .in(par_done_reg428_in),
      .write_en(par_done_reg428_write_en),
      .clk(clk),
      .out(par_done_reg428_out),
      .done(par_done_reg428_done)
  );
  
  std_reg #(1) par_done_reg429 (
      .in(par_done_reg429_in),
      .write_en(par_done_reg429_write_en),
      .clk(clk),
      .out(par_done_reg429_out),
      .done(par_done_reg429_done)
  );
  
  std_reg #(1) par_done_reg430 (
      .in(par_done_reg430_in),
      .write_en(par_done_reg430_write_en),
      .clk(clk),
      .out(par_done_reg430_out),
      .done(par_done_reg430_done)
  );
  
  std_reg #(1) par_done_reg431 (
      .in(par_done_reg431_in),
      .write_en(par_done_reg431_write_en),
      .clk(clk),
      .out(par_done_reg431_out),
      .done(par_done_reg431_done)
  );
  
  std_reg #(1) par_done_reg432 (
      .in(par_done_reg432_in),
      .write_en(par_done_reg432_write_en),
      .clk(clk),
      .out(par_done_reg432_out),
      .done(par_done_reg432_done)
  );
  
  std_reg #(1) par_done_reg433 (
      .in(par_done_reg433_in),
      .write_en(par_done_reg433_write_en),
      .clk(clk),
      .out(par_done_reg433_out),
      .done(par_done_reg433_done)
  );
  
  std_reg #(1) par_done_reg434 (
      .in(par_done_reg434_in),
      .write_en(par_done_reg434_write_en),
      .clk(clk),
      .out(par_done_reg434_out),
      .done(par_done_reg434_done)
  );
  
  std_reg #(1) par_done_reg435 (
      .in(par_done_reg435_in),
      .write_en(par_done_reg435_write_en),
      .clk(clk),
      .out(par_done_reg435_out),
      .done(par_done_reg435_done)
  );
  
  std_reg #(1) par_done_reg436 (
      .in(par_done_reg436_in),
      .write_en(par_done_reg436_write_en),
      .clk(clk),
      .out(par_done_reg436_out),
      .done(par_done_reg436_done)
  );
  
  std_reg #(1) par_done_reg437 (
      .in(par_done_reg437_in),
      .write_en(par_done_reg437_write_en),
      .clk(clk),
      .out(par_done_reg437_out),
      .done(par_done_reg437_done)
  );
  
  std_reg #(1) par_done_reg438 (
      .in(par_done_reg438_in),
      .write_en(par_done_reg438_write_en),
      .clk(clk),
      .out(par_done_reg438_out),
      .done(par_done_reg438_done)
  );
  
  std_reg #(1) par_done_reg439 (
      .in(par_done_reg439_in),
      .write_en(par_done_reg439_write_en),
      .clk(clk),
      .out(par_done_reg439_out),
      .done(par_done_reg439_done)
  );
  
  std_reg #(1) par_done_reg440 (
      .in(par_done_reg440_in),
      .write_en(par_done_reg440_write_en),
      .clk(clk),
      .out(par_done_reg440_out),
      .done(par_done_reg440_done)
  );
  
  std_reg #(1) par_done_reg441 (
      .in(par_done_reg441_in),
      .write_en(par_done_reg441_write_en),
      .clk(clk),
      .out(par_done_reg441_out),
      .done(par_done_reg441_done)
  );
  
  std_reg #(1) par_done_reg442 (
      .in(par_done_reg442_in),
      .write_en(par_done_reg442_write_en),
      .clk(clk),
      .out(par_done_reg442_out),
      .done(par_done_reg442_done)
  );
  
  std_reg #(1) par_done_reg443 (
      .in(par_done_reg443_in),
      .write_en(par_done_reg443_write_en),
      .clk(clk),
      .out(par_done_reg443_out),
      .done(par_done_reg443_done)
  );
  
  std_reg #(1) par_done_reg444 (
      .in(par_done_reg444_in),
      .write_en(par_done_reg444_write_en),
      .clk(clk),
      .out(par_done_reg444_out),
      .done(par_done_reg444_done)
  );
  
  std_reg #(1) par_done_reg445 (
      .in(par_done_reg445_in),
      .write_en(par_done_reg445_write_en),
      .clk(clk),
      .out(par_done_reg445_out),
      .done(par_done_reg445_done)
  );
  
  std_reg #(1) par_done_reg446 (
      .in(par_done_reg446_in),
      .write_en(par_done_reg446_write_en),
      .clk(clk),
      .out(par_done_reg446_out),
      .done(par_done_reg446_done)
  );
  
  std_reg #(1) par_done_reg447 (
      .in(par_done_reg447_in),
      .write_en(par_done_reg447_write_en),
      .clk(clk),
      .out(par_done_reg447_out),
      .done(par_done_reg447_done)
  );
  
  std_reg #(1) par_done_reg448 (
      .in(par_done_reg448_in),
      .write_en(par_done_reg448_write_en),
      .clk(clk),
      .out(par_done_reg448_out),
      .done(par_done_reg448_done)
  );
  
  std_reg #(1) par_done_reg449 (
      .in(par_done_reg449_in),
      .write_en(par_done_reg449_write_en),
      .clk(clk),
      .out(par_done_reg449_out),
      .done(par_done_reg449_done)
  );
  
  std_reg #(1) par_done_reg450 (
      .in(par_done_reg450_in),
      .write_en(par_done_reg450_write_en),
      .clk(clk),
      .out(par_done_reg450_out),
      .done(par_done_reg450_done)
  );
  
  std_reg #(1) par_done_reg451 (
      .in(par_done_reg451_in),
      .write_en(par_done_reg451_write_en),
      .clk(clk),
      .out(par_done_reg451_out),
      .done(par_done_reg451_done)
  );
  
  std_reg #(1) par_done_reg452 (
      .in(par_done_reg452_in),
      .write_en(par_done_reg452_write_en),
      .clk(clk),
      .out(par_done_reg452_out),
      .done(par_done_reg452_done)
  );
  
  std_reg #(1) par_done_reg453 (
      .in(par_done_reg453_in),
      .write_en(par_done_reg453_write_en),
      .clk(clk),
      .out(par_done_reg453_out),
      .done(par_done_reg453_done)
  );
  
  std_reg #(1) par_done_reg454 (
      .in(par_done_reg454_in),
      .write_en(par_done_reg454_write_en),
      .clk(clk),
      .out(par_done_reg454_out),
      .done(par_done_reg454_done)
  );
  
  std_reg #(1) par_done_reg455 (
      .in(par_done_reg455_in),
      .write_en(par_done_reg455_write_en),
      .clk(clk),
      .out(par_done_reg455_out),
      .done(par_done_reg455_done)
  );
  
  std_reg #(1) par_reset19 (
      .in(par_reset19_in),
      .write_en(par_reset19_write_en),
      .clk(clk),
      .out(par_reset19_out),
      .done(par_reset19_done)
  );
  
  std_reg #(1) par_done_reg456 (
      .in(par_done_reg456_in),
      .write_en(par_done_reg456_write_en),
      .clk(clk),
      .out(par_done_reg456_out),
      .done(par_done_reg456_done)
  );
  
  std_reg #(1) par_done_reg457 (
      .in(par_done_reg457_in),
      .write_en(par_done_reg457_write_en),
      .clk(clk),
      .out(par_done_reg457_out),
      .done(par_done_reg457_done)
  );
  
  std_reg #(1) par_done_reg458 (
      .in(par_done_reg458_in),
      .write_en(par_done_reg458_write_en),
      .clk(clk),
      .out(par_done_reg458_out),
      .done(par_done_reg458_done)
  );
  
  std_reg #(1) par_done_reg459 (
      .in(par_done_reg459_in),
      .write_en(par_done_reg459_write_en),
      .clk(clk),
      .out(par_done_reg459_out),
      .done(par_done_reg459_done)
  );
  
  std_reg #(1) par_done_reg460 (
      .in(par_done_reg460_in),
      .write_en(par_done_reg460_write_en),
      .clk(clk),
      .out(par_done_reg460_out),
      .done(par_done_reg460_done)
  );
  
  std_reg #(1) par_done_reg461 (
      .in(par_done_reg461_in),
      .write_en(par_done_reg461_write_en),
      .clk(clk),
      .out(par_done_reg461_out),
      .done(par_done_reg461_done)
  );
  
  std_reg #(1) par_done_reg462 (
      .in(par_done_reg462_in),
      .write_en(par_done_reg462_write_en),
      .clk(clk),
      .out(par_done_reg462_out),
      .done(par_done_reg462_done)
  );
  
  std_reg #(1) par_done_reg463 (
      .in(par_done_reg463_in),
      .write_en(par_done_reg463_write_en),
      .clk(clk),
      .out(par_done_reg463_out),
      .done(par_done_reg463_done)
  );
  
  std_reg #(1) par_done_reg464 (
      .in(par_done_reg464_in),
      .write_en(par_done_reg464_write_en),
      .clk(clk),
      .out(par_done_reg464_out),
      .done(par_done_reg464_done)
  );
  
  std_reg #(1) par_done_reg465 (
      .in(par_done_reg465_in),
      .write_en(par_done_reg465_write_en),
      .clk(clk),
      .out(par_done_reg465_out),
      .done(par_done_reg465_done)
  );
  
  std_reg #(1) par_done_reg466 (
      .in(par_done_reg466_in),
      .write_en(par_done_reg466_write_en),
      .clk(clk),
      .out(par_done_reg466_out),
      .done(par_done_reg466_done)
  );
  
  std_reg #(1) par_done_reg467 (
      .in(par_done_reg467_in),
      .write_en(par_done_reg467_write_en),
      .clk(clk),
      .out(par_done_reg467_out),
      .done(par_done_reg467_done)
  );
  
  std_reg #(1) par_done_reg468 (
      .in(par_done_reg468_in),
      .write_en(par_done_reg468_write_en),
      .clk(clk),
      .out(par_done_reg468_out),
      .done(par_done_reg468_done)
  );
  
  std_reg #(1) par_done_reg469 (
      .in(par_done_reg469_in),
      .write_en(par_done_reg469_write_en),
      .clk(clk),
      .out(par_done_reg469_out),
      .done(par_done_reg469_done)
  );
  
  std_reg #(1) par_done_reg470 (
      .in(par_done_reg470_in),
      .write_en(par_done_reg470_write_en),
      .clk(clk),
      .out(par_done_reg470_out),
      .done(par_done_reg470_done)
  );
  
  std_reg #(1) par_done_reg471 (
      .in(par_done_reg471_in),
      .write_en(par_done_reg471_write_en),
      .clk(clk),
      .out(par_done_reg471_out),
      .done(par_done_reg471_done)
  );
  
  std_reg #(1) par_done_reg472 (
      .in(par_done_reg472_in),
      .write_en(par_done_reg472_write_en),
      .clk(clk),
      .out(par_done_reg472_out),
      .done(par_done_reg472_done)
  );
  
  std_reg #(1) par_done_reg473 (
      .in(par_done_reg473_in),
      .write_en(par_done_reg473_write_en),
      .clk(clk),
      .out(par_done_reg473_out),
      .done(par_done_reg473_done)
  );
  
  std_reg #(1) par_done_reg474 (
      .in(par_done_reg474_in),
      .write_en(par_done_reg474_write_en),
      .clk(clk),
      .out(par_done_reg474_out),
      .done(par_done_reg474_done)
  );
  
  std_reg #(1) par_done_reg475 (
      .in(par_done_reg475_in),
      .write_en(par_done_reg475_write_en),
      .clk(clk),
      .out(par_done_reg475_out),
      .done(par_done_reg475_done)
  );
  
  std_reg #(1) par_done_reg476 (
      .in(par_done_reg476_in),
      .write_en(par_done_reg476_write_en),
      .clk(clk),
      .out(par_done_reg476_out),
      .done(par_done_reg476_done)
  );
  
  std_reg #(1) par_done_reg477 (
      .in(par_done_reg477_in),
      .write_en(par_done_reg477_write_en),
      .clk(clk),
      .out(par_done_reg477_out),
      .done(par_done_reg477_done)
  );
  
  std_reg #(1) par_done_reg478 (
      .in(par_done_reg478_in),
      .write_en(par_done_reg478_write_en),
      .clk(clk),
      .out(par_done_reg478_out),
      .done(par_done_reg478_done)
  );
  
  std_reg #(1) par_done_reg479 (
      .in(par_done_reg479_in),
      .write_en(par_done_reg479_write_en),
      .clk(clk),
      .out(par_done_reg479_out),
      .done(par_done_reg479_done)
  );
  
  std_reg #(1) par_done_reg480 (
      .in(par_done_reg480_in),
      .write_en(par_done_reg480_write_en),
      .clk(clk),
      .out(par_done_reg480_out),
      .done(par_done_reg480_done)
  );
  
  std_reg #(1) par_done_reg481 (
      .in(par_done_reg481_in),
      .write_en(par_done_reg481_write_en),
      .clk(clk),
      .out(par_done_reg481_out),
      .done(par_done_reg481_done)
  );
  
  std_reg #(1) par_done_reg482 (
      .in(par_done_reg482_in),
      .write_en(par_done_reg482_write_en),
      .clk(clk),
      .out(par_done_reg482_out),
      .done(par_done_reg482_done)
  );
  
  std_reg #(1) par_done_reg483 (
      .in(par_done_reg483_in),
      .write_en(par_done_reg483_write_en),
      .clk(clk),
      .out(par_done_reg483_out),
      .done(par_done_reg483_done)
  );
  
  std_reg #(1) par_done_reg484 (
      .in(par_done_reg484_in),
      .write_en(par_done_reg484_write_en),
      .clk(clk),
      .out(par_done_reg484_out),
      .done(par_done_reg484_done)
  );
  
  std_reg #(1) par_done_reg485 (
      .in(par_done_reg485_in),
      .write_en(par_done_reg485_write_en),
      .clk(clk),
      .out(par_done_reg485_out),
      .done(par_done_reg485_done)
  );
  
  std_reg #(1) par_done_reg486 (
      .in(par_done_reg486_in),
      .write_en(par_done_reg486_write_en),
      .clk(clk),
      .out(par_done_reg486_out),
      .done(par_done_reg486_done)
  );
  
  std_reg #(1) par_reset20 (
      .in(par_reset20_in),
      .write_en(par_reset20_write_en),
      .clk(clk),
      .out(par_reset20_out),
      .done(par_reset20_done)
  );
  
  std_reg #(1) par_done_reg487 (
      .in(par_done_reg487_in),
      .write_en(par_done_reg487_write_en),
      .clk(clk),
      .out(par_done_reg487_out),
      .done(par_done_reg487_done)
  );
  
  std_reg #(1) par_done_reg488 (
      .in(par_done_reg488_in),
      .write_en(par_done_reg488_write_en),
      .clk(clk),
      .out(par_done_reg488_out),
      .done(par_done_reg488_done)
  );
  
  std_reg #(1) par_done_reg489 (
      .in(par_done_reg489_in),
      .write_en(par_done_reg489_write_en),
      .clk(clk),
      .out(par_done_reg489_out),
      .done(par_done_reg489_done)
  );
  
  std_reg #(1) par_done_reg490 (
      .in(par_done_reg490_in),
      .write_en(par_done_reg490_write_en),
      .clk(clk),
      .out(par_done_reg490_out),
      .done(par_done_reg490_done)
  );
  
  std_reg #(1) par_done_reg491 (
      .in(par_done_reg491_in),
      .write_en(par_done_reg491_write_en),
      .clk(clk),
      .out(par_done_reg491_out),
      .done(par_done_reg491_done)
  );
  
  std_reg #(1) par_done_reg492 (
      .in(par_done_reg492_in),
      .write_en(par_done_reg492_write_en),
      .clk(clk),
      .out(par_done_reg492_out),
      .done(par_done_reg492_done)
  );
  
  std_reg #(1) par_done_reg493 (
      .in(par_done_reg493_in),
      .write_en(par_done_reg493_write_en),
      .clk(clk),
      .out(par_done_reg493_out),
      .done(par_done_reg493_done)
  );
  
  std_reg #(1) par_done_reg494 (
      .in(par_done_reg494_in),
      .write_en(par_done_reg494_write_en),
      .clk(clk),
      .out(par_done_reg494_out),
      .done(par_done_reg494_done)
  );
  
  std_reg #(1) par_done_reg495 (
      .in(par_done_reg495_in),
      .write_en(par_done_reg495_write_en),
      .clk(clk),
      .out(par_done_reg495_out),
      .done(par_done_reg495_done)
  );
  
  std_reg #(1) par_done_reg496 (
      .in(par_done_reg496_in),
      .write_en(par_done_reg496_write_en),
      .clk(clk),
      .out(par_done_reg496_out),
      .done(par_done_reg496_done)
  );
  
  std_reg #(1) par_done_reg497 (
      .in(par_done_reg497_in),
      .write_en(par_done_reg497_write_en),
      .clk(clk),
      .out(par_done_reg497_out),
      .done(par_done_reg497_done)
  );
  
  std_reg #(1) par_done_reg498 (
      .in(par_done_reg498_in),
      .write_en(par_done_reg498_write_en),
      .clk(clk),
      .out(par_done_reg498_out),
      .done(par_done_reg498_done)
  );
  
  std_reg #(1) par_done_reg499 (
      .in(par_done_reg499_in),
      .write_en(par_done_reg499_write_en),
      .clk(clk),
      .out(par_done_reg499_out),
      .done(par_done_reg499_done)
  );
  
  std_reg #(1) par_done_reg500 (
      .in(par_done_reg500_in),
      .write_en(par_done_reg500_write_en),
      .clk(clk),
      .out(par_done_reg500_out),
      .done(par_done_reg500_done)
  );
  
  std_reg #(1) par_done_reg501 (
      .in(par_done_reg501_in),
      .write_en(par_done_reg501_write_en),
      .clk(clk),
      .out(par_done_reg501_out),
      .done(par_done_reg501_done)
  );
  
  std_reg #(1) par_done_reg502 (
      .in(par_done_reg502_in),
      .write_en(par_done_reg502_write_en),
      .clk(clk),
      .out(par_done_reg502_out),
      .done(par_done_reg502_done)
  );
  
  std_reg #(1) par_done_reg503 (
      .in(par_done_reg503_in),
      .write_en(par_done_reg503_write_en),
      .clk(clk),
      .out(par_done_reg503_out),
      .done(par_done_reg503_done)
  );
  
  std_reg #(1) par_done_reg504 (
      .in(par_done_reg504_in),
      .write_en(par_done_reg504_write_en),
      .clk(clk),
      .out(par_done_reg504_out),
      .done(par_done_reg504_done)
  );
  
  std_reg #(1) par_done_reg505 (
      .in(par_done_reg505_in),
      .write_en(par_done_reg505_write_en),
      .clk(clk),
      .out(par_done_reg505_out),
      .done(par_done_reg505_done)
  );
  
  std_reg #(1) par_done_reg506 (
      .in(par_done_reg506_in),
      .write_en(par_done_reg506_write_en),
      .clk(clk),
      .out(par_done_reg506_out),
      .done(par_done_reg506_done)
  );
  
  std_reg #(1) par_done_reg507 (
      .in(par_done_reg507_in),
      .write_en(par_done_reg507_write_en),
      .clk(clk),
      .out(par_done_reg507_out),
      .done(par_done_reg507_done)
  );
  
  std_reg #(1) par_done_reg508 (
      .in(par_done_reg508_in),
      .write_en(par_done_reg508_write_en),
      .clk(clk),
      .out(par_done_reg508_out),
      .done(par_done_reg508_done)
  );
  
  std_reg #(1) par_done_reg509 (
      .in(par_done_reg509_in),
      .write_en(par_done_reg509_write_en),
      .clk(clk),
      .out(par_done_reg509_out),
      .done(par_done_reg509_done)
  );
  
  std_reg #(1) par_done_reg510 (
      .in(par_done_reg510_in),
      .write_en(par_done_reg510_write_en),
      .clk(clk),
      .out(par_done_reg510_out),
      .done(par_done_reg510_done)
  );
  
  std_reg #(1) par_done_reg511 (
      .in(par_done_reg511_in),
      .write_en(par_done_reg511_write_en),
      .clk(clk),
      .out(par_done_reg511_out),
      .done(par_done_reg511_done)
  );
  
  std_reg #(1) par_done_reg512 (
      .in(par_done_reg512_in),
      .write_en(par_done_reg512_write_en),
      .clk(clk),
      .out(par_done_reg512_out),
      .done(par_done_reg512_done)
  );
  
  std_reg #(1) par_done_reg513 (
      .in(par_done_reg513_in),
      .write_en(par_done_reg513_write_en),
      .clk(clk),
      .out(par_done_reg513_out),
      .done(par_done_reg513_done)
  );
  
  std_reg #(1) par_done_reg514 (
      .in(par_done_reg514_in),
      .write_en(par_done_reg514_write_en),
      .clk(clk),
      .out(par_done_reg514_out),
      .done(par_done_reg514_done)
  );
  
  std_reg #(1) par_done_reg515 (
      .in(par_done_reg515_in),
      .write_en(par_done_reg515_write_en),
      .clk(clk),
      .out(par_done_reg515_out),
      .done(par_done_reg515_done)
  );
  
  std_reg #(1) par_done_reg516 (
      .in(par_done_reg516_in),
      .write_en(par_done_reg516_write_en),
      .clk(clk),
      .out(par_done_reg516_out),
      .done(par_done_reg516_done)
  );
  
  std_reg #(1) par_done_reg517 (
      .in(par_done_reg517_in),
      .write_en(par_done_reg517_write_en),
      .clk(clk),
      .out(par_done_reg517_out),
      .done(par_done_reg517_done)
  );
  
  std_reg #(1) par_done_reg518 (
      .in(par_done_reg518_in),
      .write_en(par_done_reg518_write_en),
      .clk(clk),
      .out(par_done_reg518_out),
      .done(par_done_reg518_done)
  );
  
  std_reg #(1) par_done_reg519 (
      .in(par_done_reg519_in),
      .write_en(par_done_reg519_write_en),
      .clk(clk),
      .out(par_done_reg519_out),
      .done(par_done_reg519_done)
  );
  
  std_reg #(1) par_done_reg520 (
      .in(par_done_reg520_in),
      .write_en(par_done_reg520_write_en),
      .clk(clk),
      .out(par_done_reg520_out),
      .done(par_done_reg520_done)
  );
  
  std_reg #(1) par_done_reg521 (
      .in(par_done_reg521_in),
      .write_en(par_done_reg521_write_en),
      .clk(clk),
      .out(par_done_reg521_out),
      .done(par_done_reg521_done)
  );
  
  std_reg #(1) par_done_reg522 (
      .in(par_done_reg522_in),
      .write_en(par_done_reg522_write_en),
      .clk(clk),
      .out(par_done_reg522_out),
      .done(par_done_reg522_done)
  );
  
  std_reg #(1) par_done_reg523 (
      .in(par_done_reg523_in),
      .write_en(par_done_reg523_write_en),
      .clk(clk),
      .out(par_done_reg523_out),
      .done(par_done_reg523_done)
  );
  
  std_reg #(1) par_done_reg524 (
      .in(par_done_reg524_in),
      .write_en(par_done_reg524_write_en),
      .clk(clk),
      .out(par_done_reg524_out),
      .done(par_done_reg524_done)
  );
  
  std_reg #(1) par_done_reg525 (
      .in(par_done_reg525_in),
      .write_en(par_done_reg525_write_en),
      .clk(clk),
      .out(par_done_reg525_out),
      .done(par_done_reg525_done)
  );
  
  std_reg #(1) par_done_reg526 (
      .in(par_done_reg526_in),
      .write_en(par_done_reg526_write_en),
      .clk(clk),
      .out(par_done_reg526_out),
      .done(par_done_reg526_done)
  );
  
  std_reg #(1) par_done_reg527 (
      .in(par_done_reg527_in),
      .write_en(par_done_reg527_write_en),
      .clk(clk),
      .out(par_done_reg527_out),
      .done(par_done_reg527_done)
  );
  
  std_reg #(1) par_done_reg528 (
      .in(par_done_reg528_in),
      .write_en(par_done_reg528_write_en),
      .clk(clk),
      .out(par_done_reg528_out),
      .done(par_done_reg528_done)
  );
  
  std_reg #(1) par_done_reg529 (
      .in(par_done_reg529_in),
      .write_en(par_done_reg529_write_en),
      .clk(clk),
      .out(par_done_reg529_out),
      .done(par_done_reg529_done)
  );
  
  std_reg #(1) par_done_reg530 (
      .in(par_done_reg530_in),
      .write_en(par_done_reg530_write_en),
      .clk(clk),
      .out(par_done_reg530_out),
      .done(par_done_reg530_done)
  );
  
  std_reg #(1) par_done_reg531 (
      .in(par_done_reg531_in),
      .write_en(par_done_reg531_write_en),
      .clk(clk),
      .out(par_done_reg531_out),
      .done(par_done_reg531_done)
  );
  
  std_reg #(1) par_done_reg532 (
      .in(par_done_reg532_in),
      .write_en(par_done_reg532_write_en),
      .clk(clk),
      .out(par_done_reg532_out),
      .done(par_done_reg532_done)
  );
  
  std_reg #(1) par_done_reg533 (
      .in(par_done_reg533_in),
      .write_en(par_done_reg533_write_en),
      .clk(clk),
      .out(par_done_reg533_out),
      .done(par_done_reg533_done)
  );
  
  std_reg #(1) par_done_reg534 (
      .in(par_done_reg534_in),
      .write_en(par_done_reg534_write_en),
      .clk(clk),
      .out(par_done_reg534_out),
      .done(par_done_reg534_done)
  );
  
  std_reg #(1) par_done_reg535 (
      .in(par_done_reg535_in),
      .write_en(par_done_reg535_write_en),
      .clk(clk),
      .out(par_done_reg535_out),
      .done(par_done_reg535_done)
  );
  
  std_reg #(1) par_done_reg536 (
      .in(par_done_reg536_in),
      .write_en(par_done_reg536_write_en),
      .clk(clk),
      .out(par_done_reg536_out),
      .done(par_done_reg536_done)
  );
  
  std_reg #(1) par_reset21 (
      .in(par_reset21_in),
      .write_en(par_reset21_write_en),
      .clk(clk),
      .out(par_reset21_out),
      .done(par_reset21_done)
  );
  
  std_reg #(1) par_done_reg537 (
      .in(par_done_reg537_in),
      .write_en(par_done_reg537_write_en),
      .clk(clk),
      .out(par_done_reg537_out),
      .done(par_done_reg537_done)
  );
  
  std_reg #(1) par_done_reg538 (
      .in(par_done_reg538_in),
      .write_en(par_done_reg538_write_en),
      .clk(clk),
      .out(par_done_reg538_out),
      .done(par_done_reg538_done)
  );
  
  std_reg #(1) par_done_reg539 (
      .in(par_done_reg539_in),
      .write_en(par_done_reg539_write_en),
      .clk(clk),
      .out(par_done_reg539_out),
      .done(par_done_reg539_done)
  );
  
  std_reg #(1) par_done_reg540 (
      .in(par_done_reg540_in),
      .write_en(par_done_reg540_write_en),
      .clk(clk),
      .out(par_done_reg540_out),
      .done(par_done_reg540_done)
  );
  
  std_reg #(1) par_done_reg541 (
      .in(par_done_reg541_in),
      .write_en(par_done_reg541_write_en),
      .clk(clk),
      .out(par_done_reg541_out),
      .done(par_done_reg541_done)
  );
  
  std_reg #(1) par_done_reg542 (
      .in(par_done_reg542_in),
      .write_en(par_done_reg542_write_en),
      .clk(clk),
      .out(par_done_reg542_out),
      .done(par_done_reg542_done)
  );
  
  std_reg #(1) par_done_reg543 (
      .in(par_done_reg543_in),
      .write_en(par_done_reg543_write_en),
      .clk(clk),
      .out(par_done_reg543_out),
      .done(par_done_reg543_done)
  );
  
  std_reg #(1) par_done_reg544 (
      .in(par_done_reg544_in),
      .write_en(par_done_reg544_write_en),
      .clk(clk),
      .out(par_done_reg544_out),
      .done(par_done_reg544_done)
  );
  
  std_reg #(1) par_done_reg545 (
      .in(par_done_reg545_in),
      .write_en(par_done_reg545_write_en),
      .clk(clk),
      .out(par_done_reg545_out),
      .done(par_done_reg545_done)
  );
  
  std_reg #(1) par_done_reg546 (
      .in(par_done_reg546_in),
      .write_en(par_done_reg546_write_en),
      .clk(clk),
      .out(par_done_reg546_out),
      .done(par_done_reg546_done)
  );
  
  std_reg #(1) par_done_reg547 (
      .in(par_done_reg547_in),
      .write_en(par_done_reg547_write_en),
      .clk(clk),
      .out(par_done_reg547_out),
      .done(par_done_reg547_done)
  );
  
  std_reg #(1) par_done_reg548 (
      .in(par_done_reg548_in),
      .write_en(par_done_reg548_write_en),
      .clk(clk),
      .out(par_done_reg548_out),
      .done(par_done_reg548_done)
  );
  
  std_reg #(1) par_done_reg549 (
      .in(par_done_reg549_in),
      .write_en(par_done_reg549_write_en),
      .clk(clk),
      .out(par_done_reg549_out),
      .done(par_done_reg549_done)
  );
  
  std_reg #(1) par_done_reg550 (
      .in(par_done_reg550_in),
      .write_en(par_done_reg550_write_en),
      .clk(clk),
      .out(par_done_reg550_out),
      .done(par_done_reg550_done)
  );
  
  std_reg #(1) par_done_reg551 (
      .in(par_done_reg551_in),
      .write_en(par_done_reg551_write_en),
      .clk(clk),
      .out(par_done_reg551_out),
      .done(par_done_reg551_done)
  );
  
  std_reg #(1) par_done_reg552 (
      .in(par_done_reg552_in),
      .write_en(par_done_reg552_write_en),
      .clk(clk),
      .out(par_done_reg552_out),
      .done(par_done_reg552_done)
  );
  
  std_reg #(1) par_done_reg553 (
      .in(par_done_reg553_in),
      .write_en(par_done_reg553_write_en),
      .clk(clk),
      .out(par_done_reg553_out),
      .done(par_done_reg553_done)
  );
  
  std_reg #(1) par_done_reg554 (
      .in(par_done_reg554_in),
      .write_en(par_done_reg554_write_en),
      .clk(clk),
      .out(par_done_reg554_out),
      .done(par_done_reg554_done)
  );
  
  std_reg #(1) par_done_reg555 (
      .in(par_done_reg555_in),
      .write_en(par_done_reg555_write_en),
      .clk(clk),
      .out(par_done_reg555_out),
      .done(par_done_reg555_done)
  );
  
  std_reg #(1) par_done_reg556 (
      .in(par_done_reg556_in),
      .write_en(par_done_reg556_write_en),
      .clk(clk),
      .out(par_done_reg556_out),
      .done(par_done_reg556_done)
  );
  
  std_reg #(1) par_done_reg557 (
      .in(par_done_reg557_in),
      .write_en(par_done_reg557_write_en),
      .clk(clk),
      .out(par_done_reg557_out),
      .done(par_done_reg557_done)
  );
  
  std_reg #(1) par_done_reg558 (
      .in(par_done_reg558_in),
      .write_en(par_done_reg558_write_en),
      .clk(clk),
      .out(par_done_reg558_out),
      .done(par_done_reg558_done)
  );
  
  std_reg #(1) par_done_reg559 (
      .in(par_done_reg559_in),
      .write_en(par_done_reg559_write_en),
      .clk(clk),
      .out(par_done_reg559_out),
      .done(par_done_reg559_done)
  );
  
  std_reg #(1) par_done_reg560 (
      .in(par_done_reg560_in),
      .write_en(par_done_reg560_write_en),
      .clk(clk),
      .out(par_done_reg560_out),
      .done(par_done_reg560_done)
  );
  
  std_reg #(1) par_done_reg561 (
      .in(par_done_reg561_in),
      .write_en(par_done_reg561_write_en),
      .clk(clk),
      .out(par_done_reg561_out),
      .done(par_done_reg561_done)
  );
  
  std_reg #(1) par_done_reg562 (
      .in(par_done_reg562_in),
      .write_en(par_done_reg562_write_en),
      .clk(clk),
      .out(par_done_reg562_out),
      .done(par_done_reg562_done)
  );
  
  std_reg #(1) par_done_reg563 (
      .in(par_done_reg563_in),
      .write_en(par_done_reg563_write_en),
      .clk(clk),
      .out(par_done_reg563_out),
      .done(par_done_reg563_done)
  );
  
  std_reg #(1) par_reset22 (
      .in(par_reset22_in),
      .write_en(par_reset22_write_en),
      .clk(clk),
      .out(par_reset22_out),
      .done(par_reset22_done)
  );
  
  std_reg #(1) par_done_reg564 (
      .in(par_done_reg564_in),
      .write_en(par_done_reg564_write_en),
      .clk(clk),
      .out(par_done_reg564_out),
      .done(par_done_reg564_done)
  );
  
  std_reg #(1) par_done_reg565 (
      .in(par_done_reg565_in),
      .write_en(par_done_reg565_write_en),
      .clk(clk),
      .out(par_done_reg565_out),
      .done(par_done_reg565_done)
  );
  
  std_reg #(1) par_done_reg566 (
      .in(par_done_reg566_in),
      .write_en(par_done_reg566_write_en),
      .clk(clk),
      .out(par_done_reg566_out),
      .done(par_done_reg566_done)
  );
  
  std_reg #(1) par_done_reg567 (
      .in(par_done_reg567_in),
      .write_en(par_done_reg567_write_en),
      .clk(clk),
      .out(par_done_reg567_out),
      .done(par_done_reg567_done)
  );
  
  std_reg #(1) par_done_reg568 (
      .in(par_done_reg568_in),
      .write_en(par_done_reg568_write_en),
      .clk(clk),
      .out(par_done_reg568_out),
      .done(par_done_reg568_done)
  );
  
  std_reg #(1) par_done_reg569 (
      .in(par_done_reg569_in),
      .write_en(par_done_reg569_write_en),
      .clk(clk),
      .out(par_done_reg569_out),
      .done(par_done_reg569_done)
  );
  
  std_reg #(1) par_done_reg570 (
      .in(par_done_reg570_in),
      .write_en(par_done_reg570_write_en),
      .clk(clk),
      .out(par_done_reg570_out),
      .done(par_done_reg570_done)
  );
  
  std_reg #(1) par_done_reg571 (
      .in(par_done_reg571_in),
      .write_en(par_done_reg571_write_en),
      .clk(clk),
      .out(par_done_reg571_out),
      .done(par_done_reg571_done)
  );
  
  std_reg #(1) par_done_reg572 (
      .in(par_done_reg572_in),
      .write_en(par_done_reg572_write_en),
      .clk(clk),
      .out(par_done_reg572_out),
      .done(par_done_reg572_done)
  );
  
  std_reg #(1) par_done_reg573 (
      .in(par_done_reg573_in),
      .write_en(par_done_reg573_write_en),
      .clk(clk),
      .out(par_done_reg573_out),
      .done(par_done_reg573_done)
  );
  
  std_reg #(1) par_done_reg574 (
      .in(par_done_reg574_in),
      .write_en(par_done_reg574_write_en),
      .clk(clk),
      .out(par_done_reg574_out),
      .done(par_done_reg574_done)
  );
  
  std_reg #(1) par_done_reg575 (
      .in(par_done_reg575_in),
      .write_en(par_done_reg575_write_en),
      .clk(clk),
      .out(par_done_reg575_out),
      .done(par_done_reg575_done)
  );
  
  std_reg #(1) par_done_reg576 (
      .in(par_done_reg576_in),
      .write_en(par_done_reg576_write_en),
      .clk(clk),
      .out(par_done_reg576_out),
      .done(par_done_reg576_done)
  );
  
  std_reg #(1) par_done_reg577 (
      .in(par_done_reg577_in),
      .write_en(par_done_reg577_write_en),
      .clk(clk),
      .out(par_done_reg577_out),
      .done(par_done_reg577_done)
  );
  
  std_reg #(1) par_done_reg578 (
      .in(par_done_reg578_in),
      .write_en(par_done_reg578_write_en),
      .clk(clk),
      .out(par_done_reg578_out),
      .done(par_done_reg578_done)
  );
  
  std_reg #(1) par_done_reg579 (
      .in(par_done_reg579_in),
      .write_en(par_done_reg579_write_en),
      .clk(clk),
      .out(par_done_reg579_out),
      .done(par_done_reg579_done)
  );
  
  std_reg #(1) par_done_reg580 (
      .in(par_done_reg580_in),
      .write_en(par_done_reg580_write_en),
      .clk(clk),
      .out(par_done_reg580_out),
      .done(par_done_reg580_done)
  );
  
  std_reg #(1) par_done_reg581 (
      .in(par_done_reg581_in),
      .write_en(par_done_reg581_write_en),
      .clk(clk),
      .out(par_done_reg581_out),
      .done(par_done_reg581_done)
  );
  
  std_reg #(1) par_done_reg582 (
      .in(par_done_reg582_in),
      .write_en(par_done_reg582_write_en),
      .clk(clk),
      .out(par_done_reg582_out),
      .done(par_done_reg582_done)
  );
  
  std_reg #(1) par_done_reg583 (
      .in(par_done_reg583_in),
      .write_en(par_done_reg583_write_en),
      .clk(clk),
      .out(par_done_reg583_out),
      .done(par_done_reg583_done)
  );
  
  std_reg #(1) par_done_reg584 (
      .in(par_done_reg584_in),
      .write_en(par_done_reg584_write_en),
      .clk(clk),
      .out(par_done_reg584_out),
      .done(par_done_reg584_done)
  );
  
  std_reg #(1) par_done_reg585 (
      .in(par_done_reg585_in),
      .write_en(par_done_reg585_write_en),
      .clk(clk),
      .out(par_done_reg585_out),
      .done(par_done_reg585_done)
  );
  
  std_reg #(1) par_done_reg586 (
      .in(par_done_reg586_in),
      .write_en(par_done_reg586_write_en),
      .clk(clk),
      .out(par_done_reg586_out),
      .done(par_done_reg586_done)
  );
  
  std_reg #(1) par_done_reg587 (
      .in(par_done_reg587_in),
      .write_en(par_done_reg587_write_en),
      .clk(clk),
      .out(par_done_reg587_out),
      .done(par_done_reg587_done)
  );
  
  std_reg #(1) par_done_reg588 (
      .in(par_done_reg588_in),
      .write_en(par_done_reg588_write_en),
      .clk(clk),
      .out(par_done_reg588_out),
      .done(par_done_reg588_done)
  );
  
  std_reg #(1) par_done_reg589 (
      .in(par_done_reg589_in),
      .write_en(par_done_reg589_write_en),
      .clk(clk),
      .out(par_done_reg589_out),
      .done(par_done_reg589_done)
  );
  
  std_reg #(1) par_done_reg590 (
      .in(par_done_reg590_in),
      .write_en(par_done_reg590_write_en),
      .clk(clk),
      .out(par_done_reg590_out),
      .done(par_done_reg590_done)
  );
  
  std_reg #(1) par_done_reg591 (
      .in(par_done_reg591_in),
      .write_en(par_done_reg591_write_en),
      .clk(clk),
      .out(par_done_reg591_out),
      .done(par_done_reg591_done)
  );
  
  std_reg #(1) par_done_reg592 (
      .in(par_done_reg592_in),
      .write_en(par_done_reg592_write_en),
      .clk(clk),
      .out(par_done_reg592_out),
      .done(par_done_reg592_done)
  );
  
  std_reg #(1) par_done_reg593 (
      .in(par_done_reg593_in),
      .write_en(par_done_reg593_write_en),
      .clk(clk),
      .out(par_done_reg593_out),
      .done(par_done_reg593_done)
  );
  
  std_reg #(1) par_done_reg594 (
      .in(par_done_reg594_in),
      .write_en(par_done_reg594_write_en),
      .clk(clk),
      .out(par_done_reg594_out),
      .done(par_done_reg594_done)
  );
  
  std_reg #(1) par_done_reg595 (
      .in(par_done_reg595_in),
      .write_en(par_done_reg595_write_en),
      .clk(clk),
      .out(par_done_reg595_out),
      .done(par_done_reg595_done)
  );
  
  std_reg #(1) par_done_reg596 (
      .in(par_done_reg596_in),
      .write_en(par_done_reg596_write_en),
      .clk(clk),
      .out(par_done_reg596_out),
      .done(par_done_reg596_done)
  );
  
  std_reg #(1) par_done_reg597 (
      .in(par_done_reg597_in),
      .write_en(par_done_reg597_write_en),
      .clk(clk),
      .out(par_done_reg597_out),
      .done(par_done_reg597_done)
  );
  
  std_reg #(1) par_done_reg598 (
      .in(par_done_reg598_in),
      .write_en(par_done_reg598_write_en),
      .clk(clk),
      .out(par_done_reg598_out),
      .done(par_done_reg598_done)
  );
  
  std_reg #(1) par_done_reg599 (
      .in(par_done_reg599_in),
      .write_en(par_done_reg599_write_en),
      .clk(clk),
      .out(par_done_reg599_out),
      .done(par_done_reg599_done)
  );
  
  std_reg #(1) par_done_reg600 (
      .in(par_done_reg600_in),
      .write_en(par_done_reg600_write_en),
      .clk(clk),
      .out(par_done_reg600_out),
      .done(par_done_reg600_done)
  );
  
  std_reg #(1) par_done_reg601 (
      .in(par_done_reg601_in),
      .write_en(par_done_reg601_write_en),
      .clk(clk),
      .out(par_done_reg601_out),
      .done(par_done_reg601_done)
  );
  
  std_reg #(1) par_done_reg602 (
      .in(par_done_reg602_in),
      .write_en(par_done_reg602_write_en),
      .clk(clk),
      .out(par_done_reg602_out),
      .done(par_done_reg602_done)
  );
  
  std_reg #(1) par_done_reg603 (
      .in(par_done_reg603_in),
      .write_en(par_done_reg603_write_en),
      .clk(clk),
      .out(par_done_reg603_out),
      .done(par_done_reg603_done)
  );
  
  std_reg #(1) par_done_reg604 (
      .in(par_done_reg604_in),
      .write_en(par_done_reg604_write_en),
      .clk(clk),
      .out(par_done_reg604_out),
      .done(par_done_reg604_done)
  );
  
  std_reg #(1) par_done_reg605 (
      .in(par_done_reg605_in),
      .write_en(par_done_reg605_write_en),
      .clk(clk),
      .out(par_done_reg605_out),
      .done(par_done_reg605_done)
  );
  
  std_reg #(1) par_reset23 (
      .in(par_reset23_in),
      .write_en(par_reset23_write_en),
      .clk(clk),
      .out(par_reset23_out),
      .done(par_reset23_done)
  );
  
  std_reg #(1) par_done_reg606 (
      .in(par_done_reg606_in),
      .write_en(par_done_reg606_write_en),
      .clk(clk),
      .out(par_done_reg606_out),
      .done(par_done_reg606_done)
  );
  
  std_reg #(1) par_done_reg607 (
      .in(par_done_reg607_in),
      .write_en(par_done_reg607_write_en),
      .clk(clk),
      .out(par_done_reg607_out),
      .done(par_done_reg607_done)
  );
  
  std_reg #(1) par_done_reg608 (
      .in(par_done_reg608_in),
      .write_en(par_done_reg608_write_en),
      .clk(clk),
      .out(par_done_reg608_out),
      .done(par_done_reg608_done)
  );
  
  std_reg #(1) par_done_reg609 (
      .in(par_done_reg609_in),
      .write_en(par_done_reg609_write_en),
      .clk(clk),
      .out(par_done_reg609_out),
      .done(par_done_reg609_done)
  );
  
  std_reg #(1) par_done_reg610 (
      .in(par_done_reg610_in),
      .write_en(par_done_reg610_write_en),
      .clk(clk),
      .out(par_done_reg610_out),
      .done(par_done_reg610_done)
  );
  
  std_reg #(1) par_done_reg611 (
      .in(par_done_reg611_in),
      .write_en(par_done_reg611_write_en),
      .clk(clk),
      .out(par_done_reg611_out),
      .done(par_done_reg611_done)
  );
  
  std_reg #(1) par_done_reg612 (
      .in(par_done_reg612_in),
      .write_en(par_done_reg612_write_en),
      .clk(clk),
      .out(par_done_reg612_out),
      .done(par_done_reg612_done)
  );
  
  std_reg #(1) par_done_reg613 (
      .in(par_done_reg613_in),
      .write_en(par_done_reg613_write_en),
      .clk(clk),
      .out(par_done_reg613_out),
      .done(par_done_reg613_done)
  );
  
  std_reg #(1) par_done_reg614 (
      .in(par_done_reg614_in),
      .write_en(par_done_reg614_write_en),
      .clk(clk),
      .out(par_done_reg614_out),
      .done(par_done_reg614_done)
  );
  
  std_reg #(1) par_done_reg615 (
      .in(par_done_reg615_in),
      .write_en(par_done_reg615_write_en),
      .clk(clk),
      .out(par_done_reg615_out),
      .done(par_done_reg615_done)
  );
  
  std_reg #(1) par_done_reg616 (
      .in(par_done_reg616_in),
      .write_en(par_done_reg616_write_en),
      .clk(clk),
      .out(par_done_reg616_out),
      .done(par_done_reg616_done)
  );
  
  std_reg #(1) par_done_reg617 (
      .in(par_done_reg617_in),
      .write_en(par_done_reg617_write_en),
      .clk(clk),
      .out(par_done_reg617_out),
      .done(par_done_reg617_done)
  );
  
  std_reg #(1) par_done_reg618 (
      .in(par_done_reg618_in),
      .write_en(par_done_reg618_write_en),
      .clk(clk),
      .out(par_done_reg618_out),
      .done(par_done_reg618_done)
  );
  
  std_reg #(1) par_done_reg619 (
      .in(par_done_reg619_in),
      .write_en(par_done_reg619_write_en),
      .clk(clk),
      .out(par_done_reg619_out),
      .done(par_done_reg619_done)
  );
  
  std_reg #(1) par_done_reg620 (
      .in(par_done_reg620_in),
      .write_en(par_done_reg620_write_en),
      .clk(clk),
      .out(par_done_reg620_out),
      .done(par_done_reg620_done)
  );
  
  std_reg #(1) par_done_reg621 (
      .in(par_done_reg621_in),
      .write_en(par_done_reg621_write_en),
      .clk(clk),
      .out(par_done_reg621_out),
      .done(par_done_reg621_done)
  );
  
  std_reg #(1) par_done_reg622 (
      .in(par_done_reg622_in),
      .write_en(par_done_reg622_write_en),
      .clk(clk),
      .out(par_done_reg622_out),
      .done(par_done_reg622_done)
  );
  
  std_reg #(1) par_done_reg623 (
      .in(par_done_reg623_in),
      .write_en(par_done_reg623_write_en),
      .clk(clk),
      .out(par_done_reg623_out),
      .done(par_done_reg623_done)
  );
  
  std_reg #(1) par_done_reg624 (
      .in(par_done_reg624_in),
      .write_en(par_done_reg624_write_en),
      .clk(clk),
      .out(par_done_reg624_out),
      .done(par_done_reg624_done)
  );
  
  std_reg #(1) par_done_reg625 (
      .in(par_done_reg625_in),
      .write_en(par_done_reg625_write_en),
      .clk(clk),
      .out(par_done_reg625_out),
      .done(par_done_reg625_done)
  );
  
  std_reg #(1) par_done_reg626 (
      .in(par_done_reg626_in),
      .write_en(par_done_reg626_write_en),
      .clk(clk),
      .out(par_done_reg626_out),
      .done(par_done_reg626_done)
  );
  
  std_reg #(1) par_reset24 (
      .in(par_reset24_in),
      .write_en(par_reset24_write_en),
      .clk(clk),
      .out(par_reset24_out),
      .done(par_reset24_done)
  );
  
  std_reg #(1) par_done_reg627 (
      .in(par_done_reg627_in),
      .write_en(par_done_reg627_write_en),
      .clk(clk),
      .out(par_done_reg627_out),
      .done(par_done_reg627_done)
  );
  
  std_reg #(1) par_done_reg628 (
      .in(par_done_reg628_in),
      .write_en(par_done_reg628_write_en),
      .clk(clk),
      .out(par_done_reg628_out),
      .done(par_done_reg628_done)
  );
  
  std_reg #(1) par_done_reg629 (
      .in(par_done_reg629_in),
      .write_en(par_done_reg629_write_en),
      .clk(clk),
      .out(par_done_reg629_out),
      .done(par_done_reg629_done)
  );
  
  std_reg #(1) par_done_reg630 (
      .in(par_done_reg630_in),
      .write_en(par_done_reg630_write_en),
      .clk(clk),
      .out(par_done_reg630_out),
      .done(par_done_reg630_done)
  );
  
  std_reg #(1) par_done_reg631 (
      .in(par_done_reg631_in),
      .write_en(par_done_reg631_write_en),
      .clk(clk),
      .out(par_done_reg631_out),
      .done(par_done_reg631_done)
  );
  
  std_reg #(1) par_done_reg632 (
      .in(par_done_reg632_in),
      .write_en(par_done_reg632_write_en),
      .clk(clk),
      .out(par_done_reg632_out),
      .done(par_done_reg632_done)
  );
  
  std_reg #(1) par_done_reg633 (
      .in(par_done_reg633_in),
      .write_en(par_done_reg633_write_en),
      .clk(clk),
      .out(par_done_reg633_out),
      .done(par_done_reg633_done)
  );
  
  std_reg #(1) par_done_reg634 (
      .in(par_done_reg634_in),
      .write_en(par_done_reg634_write_en),
      .clk(clk),
      .out(par_done_reg634_out),
      .done(par_done_reg634_done)
  );
  
  std_reg #(1) par_done_reg635 (
      .in(par_done_reg635_in),
      .write_en(par_done_reg635_write_en),
      .clk(clk),
      .out(par_done_reg635_out),
      .done(par_done_reg635_done)
  );
  
  std_reg #(1) par_done_reg636 (
      .in(par_done_reg636_in),
      .write_en(par_done_reg636_write_en),
      .clk(clk),
      .out(par_done_reg636_out),
      .done(par_done_reg636_done)
  );
  
  std_reg #(1) par_done_reg637 (
      .in(par_done_reg637_in),
      .write_en(par_done_reg637_write_en),
      .clk(clk),
      .out(par_done_reg637_out),
      .done(par_done_reg637_done)
  );
  
  std_reg #(1) par_done_reg638 (
      .in(par_done_reg638_in),
      .write_en(par_done_reg638_write_en),
      .clk(clk),
      .out(par_done_reg638_out),
      .done(par_done_reg638_done)
  );
  
  std_reg #(1) par_done_reg639 (
      .in(par_done_reg639_in),
      .write_en(par_done_reg639_write_en),
      .clk(clk),
      .out(par_done_reg639_out),
      .done(par_done_reg639_done)
  );
  
  std_reg #(1) par_done_reg640 (
      .in(par_done_reg640_in),
      .write_en(par_done_reg640_write_en),
      .clk(clk),
      .out(par_done_reg640_out),
      .done(par_done_reg640_done)
  );
  
  std_reg #(1) par_done_reg641 (
      .in(par_done_reg641_in),
      .write_en(par_done_reg641_write_en),
      .clk(clk),
      .out(par_done_reg641_out),
      .done(par_done_reg641_done)
  );
  
  std_reg #(1) par_done_reg642 (
      .in(par_done_reg642_in),
      .write_en(par_done_reg642_write_en),
      .clk(clk),
      .out(par_done_reg642_out),
      .done(par_done_reg642_done)
  );
  
  std_reg #(1) par_done_reg643 (
      .in(par_done_reg643_in),
      .write_en(par_done_reg643_write_en),
      .clk(clk),
      .out(par_done_reg643_out),
      .done(par_done_reg643_done)
  );
  
  std_reg #(1) par_done_reg644 (
      .in(par_done_reg644_in),
      .write_en(par_done_reg644_write_en),
      .clk(clk),
      .out(par_done_reg644_out),
      .done(par_done_reg644_done)
  );
  
  std_reg #(1) par_done_reg645 (
      .in(par_done_reg645_in),
      .write_en(par_done_reg645_write_en),
      .clk(clk),
      .out(par_done_reg645_out),
      .done(par_done_reg645_done)
  );
  
  std_reg #(1) par_done_reg646 (
      .in(par_done_reg646_in),
      .write_en(par_done_reg646_write_en),
      .clk(clk),
      .out(par_done_reg646_out),
      .done(par_done_reg646_done)
  );
  
  std_reg #(1) par_done_reg647 (
      .in(par_done_reg647_in),
      .write_en(par_done_reg647_write_en),
      .clk(clk),
      .out(par_done_reg647_out),
      .done(par_done_reg647_done)
  );
  
  std_reg #(1) par_done_reg648 (
      .in(par_done_reg648_in),
      .write_en(par_done_reg648_write_en),
      .clk(clk),
      .out(par_done_reg648_out),
      .done(par_done_reg648_done)
  );
  
  std_reg #(1) par_done_reg649 (
      .in(par_done_reg649_in),
      .write_en(par_done_reg649_write_en),
      .clk(clk),
      .out(par_done_reg649_out),
      .done(par_done_reg649_done)
  );
  
  std_reg #(1) par_done_reg650 (
      .in(par_done_reg650_in),
      .write_en(par_done_reg650_write_en),
      .clk(clk),
      .out(par_done_reg650_out),
      .done(par_done_reg650_done)
  );
  
  std_reg #(1) par_done_reg651 (
      .in(par_done_reg651_in),
      .write_en(par_done_reg651_write_en),
      .clk(clk),
      .out(par_done_reg651_out),
      .done(par_done_reg651_done)
  );
  
  std_reg #(1) par_done_reg652 (
      .in(par_done_reg652_in),
      .write_en(par_done_reg652_write_en),
      .clk(clk),
      .out(par_done_reg652_out),
      .done(par_done_reg652_done)
  );
  
  std_reg #(1) par_done_reg653 (
      .in(par_done_reg653_in),
      .write_en(par_done_reg653_write_en),
      .clk(clk),
      .out(par_done_reg653_out),
      .done(par_done_reg653_done)
  );
  
  std_reg #(1) par_done_reg654 (
      .in(par_done_reg654_in),
      .write_en(par_done_reg654_write_en),
      .clk(clk),
      .out(par_done_reg654_out),
      .done(par_done_reg654_done)
  );
  
  std_reg #(1) par_done_reg655 (
      .in(par_done_reg655_in),
      .write_en(par_done_reg655_write_en),
      .clk(clk),
      .out(par_done_reg655_out),
      .done(par_done_reg655_done)
  );
  
  std_reg #(1) par_done_reg656 (
      .in(par_done_reg656_in),
      .write_en(par_done_reg656_write_en),
      .clk(clk),
      .out(par_done_reg656_out),
      .done(par_done_reg656_done)
  );
  
  std_reg #(1) par_reset25 (
      .in(par_reset25_in),
      .write_en(par_reset25_write_en),
      .clk(clk),
      .out(par_reset25_out),
      .done(par_reset25_done)
  );
  
  std_reg #(1) par_done_reg657 (
      .in(par_done_reg657_in),
      .write_en(par_done_reg657_write_en),
      .clk(clk),
      .out(par_done_reg657_out),
      .done(par_done_reg657_done)
  );
  
  std_reg #(1) par_done_reg658 (
      .in(par_done_reg658_in),
      .write_en(par_done_reg658_write_en),
      .clk(clk),
      .out(par_done_reg658_out),
      .done(par_done_reg658_done)
  );
  
  std_reg #(1) par_done_reg659 (
      .in(par_done_reg659_in),
      .write_en(par_done_reg659_write_en),
      .clk(clk),
      .out(par_done_reg659_out),
      .done(par_done_reg659_done)
  );
  
  std_reg #(1) par_done_reg660 (
      .in(par_done_reg660_in),
      .write_en(par_done_reg660_write_en),
      .clk(clk),
      .out(par_done_reg660_out),
      .done(par_done_reg660_done)
  );
  
  std_reg #(1) par_done_reg661 (
      .in(par_done_reg661_in),
      .write_en(par_done_reg661_write_en),
      .clk(clk),
      .out(par_done_reg661_out),
      .done(par_done_reg661_done)
  );
  
  std_reg #(1) par_done_reg662 (
      .in(par_done_reg662_in),
      .write_en(par_done_reg662_write_en),
      .clk(clk),
      .out(par_done_reg662_out),
      .done(par_done_reg662_done)
  );
  
  std_reg #(1) par_done_reg663 (
      .in(par_done_reg663_in),
      .write_en(par_done_reg663_write_en),
      .clk(clk),
      .out(par_done_reg663_out),
      .done(par_done_reg663_done)
  );
  
  std_reg #(1) par_done_reg664 (
      .in(par_done_reg664_in),
      .write_en(par_done_reg664_write_en),
      .clk(clk),
      .out(par_done_reg664_out),
      .done(par_done_reg664_done)
  );
  
  std_reg #(1) par_done_reg665 (
      .in(par_done_reg665_in),
      .write_en(par_done_reg665_write_en),
      .clk(clk),
      .out(par_done_reg665_out),
      .done(par_done_reg665_done)
  );
  
  std_reg #(1) par_done_reg666 (
      .in(par_done_reg666_in),
      .write_en(par_done_reg666_write_en),
      .clk(clk),
      .out(par_done_reg666_out),
      .done(par_done_reg666_done)
  );
  
  std_reg #(1) par_done_reg667 (
      .in(par_done_reg667_in),
      .write_en(par_done_reg667_write_en),
      .clk(clk),
      .out(par_done_reg667_out),
      .done(par_done_reg667_done)
  );
  
  std_reg #(1) par_done_reg668 (
      .in(par_done_reg668_in),
      .write_en(par_done_reg668_write_en),
      .clk(clk),
      .out(par_done_reg668_out),
      .done(par_done_reg668_done)
  );
  
  std_reg #(1) par_done_reg669 (
      .in(par_done_reg669_in),
      .write_en(par_done_reg669_write_en),
      .clk(clk),
      .out(par_done_reg669_out),
      .done(par_done_reg669_done)
  );
  
  std_reg #(1) par_done_reg670 (
      .in(par_done_reg670_in),
      .write_en(par_done_reg670_write_en),
      .clk(clk),
      .out(par_done_reg670_out),
      .done(par_done_reg670_done)
  );
  
  std_reg #(1) par_done_reg671 (
      .in(par_done_reg671_in),
      .write_en(par_done_reg671_write_en),
      .clk(clk),
      .out(par_done_reg671_out),
      .done(par_done_reg671_done)
  );
  
  std_reg #(1) par_reset26 (
      .in(par_reset26_in),
      .write_en(par_reset26_write_en),
      .clk(clk),
      .out(par_reset26_out),
      .done(par_reset26_done)
  );
  
  std_reg #(1) par_done_reg672 (
      .in(par_done_reg672_in),
      .write_en(par_done_reg672_write_en),
      .clk(clk),
      .out(par_done_reg672_out),
      .done(par_done_reg672_done)
  );
  
  std_reg #(1) par_done_reg673 (
      .in(par_done_reg673_in),
      .write_en(par_done_reg673_write_en),
      .clk(clk),
      .out(par_done_reg673_out),
      .done(par_done_reg673_done)
  );
  
  std_reg #(1) par_done_reg674 (
      .in(par_done_reg674_in),
      .write_en(par_done_reg674_write_en),
      .clk(clk),
      .out(par_done_reg674_out),
      .done(par_done_reg674_done)
  );
  
  std_reg #(1) par_done_reg675 (
      .in(par_done_reg675_in),
      .write_en(par_done_reg675_write_en),
      .clk(clk),
      .out(par_done_reg675_out),
      .done(par_done_reg675_done)
  );
  
  std_reg #(1) par_done_reg676 (
      .in(par_done_reg676_in),
      .write_en(par_done_reg676_write_en),
      .clk(clk),
      .out(par_done_reg676_out),
      .done(par_done_reg676_done)
  );
  
  std_reg #(1) par_done_reg677 (
      .in(par_done_reg677_in),
      .write_en(par_done_reg677_write_en),
      .clk(clk),
      .out(par_done_reg677_out),
      .done(par_done_reg677_done)
  );
  
  std_reg #(1) par_done_reg678 (
      .in(par_done_reg678_in),
      .write_en(par_done_reg678_write_en),
      .clk(clk),
      .out(par_done_reg678_out),
      .done(par_done_reg678_done)
  );
  
  std_reg #(1) par_done_reg679 (
      .in(par_done_reg679_in),
      .write_en(par_done_reg679_write_en),
      .clk(clk),
      .out(par_done_reg679_out),
      .done(par_done_reg679_done)
  );
  
  std_reg #(1) par_done_reg680 (
      .in(par_done_reg680_in),
      .write_en(par_done_reg680_write_en),
      .clk(clk),
      .out(par_done_reg680_out),
      .done(par_done_reg680_done)
  );
  
  std_reg #(1) par_done_reg681 (
      .in(par_done_reg681_in),
      .write_en(par_done_reg681_write_en),
      .clk(clk),
      .out(par_done_reg681_out),
      .done(par_done_reg681_done)
  );
  
  std_reg #(1) par_done_reg682 (
      .in(par_done_reg682_in),
      .write_en(par_done_reg682_write_en),
      .clk(clk),
      .out(par_done_reg682_out),
      .done(par_done_reg682_done)
  );
  
  std_reg #(1) par_done_reg683 (
      .in(par_done_reg683_in),
      .write_en(par_done_reg683_write_en),
      .clk(clk),
      .out(par_done_reg683_out),
      .done(par_done_reg683_done)
  );
  
  std_reg #(1) par_done_reg684 (
      .in(par_done_reg684_in),
      .write_en(par_done_reg684_write_en),
      .clk(clk),
      .out(par_done_reg684_out),
      .done(par_done_reg684_done)
  );
  
  std_reg #(1) par_done_reg685 (
      .in(par_done_reg685_in),
      .write_en(par_done_reg685_write_en),
      .clk(clk),
      .out(par_done_reg685_out),
      .done(par_done_reg685_done)
  );
  
  std_reg #(1) par_done_reg686 (
      .in(par_done_reg686_in),
      .write_en(par_done_reg686_write_en),
      .clk(clk),
      .out(par_done_reg686_out),
      .done(par_done_reg686_done)
  );
  
  std_reg #(1) par_done_reg687 (
      .in(par_done_reg687_in),
      .write_en(par_done_reg687_write_en),
      .clk(clk),
      .out(par_done_reg687_out),
      .done(par_done_reg687_done)
  );
  
  std_reg #(1) par_done_reg688 (
      .in(par_done_reg688_in),
      .write_en(par_done_reg688_write_en),
      .clk(clk),
      .out(par_done_reg688_out),
      .done(par_done_reg688_done)
  );
  
  std_reg #(1) par_done_reg689 (
      .in(par_done_reg689_in),
      .write_en(par_done_reg689_write_en),
      .clk(clk),
      .out(par_done_reg689_out),
      .done(par_done_reg689_done)
  );
  
  std_reg #(1) par_done_reg690 (
      .in(par_done_reg690_in),
      .write_en(par_done_reg690_write_en),
      .clk(clk),
      .out(par_done_reg690_out),
      .done(par_done_reg690_done)
  );
  
  std_reg #(1) par_done_reg691 (
      .in(par_done_reg691_in),
      .write_en(par_done_reg691_write_en),
      .clk(clk),
      .out(par_done_reg691_out),
      .done(par_done_reg691_done)
  );
  
  std_reg #(1) par_reset27 (
      .in(par_reset27_in),
      .write_en(par_reset27_write_en),
      .clk(clk),
      .out(par_reset27_out),
      .done(par_reset27_done)
  );
  
  std_reg #(1) par_done_reg692 (
      .in(par_done_reg692_in),
      .write_en(par_done_reg692_write_en),
      .clk(clk),
      .out(par_done_reg692_out),
      .done(par_done_reg692_done)
  );
  
  std_reg #(1) par_done_reg693 (
      .in(par_done_reg693_in),
      .write_en(par_done_reg693_write_en),
      .clk(clk),
      .out(par_done_reg693_out),
      .done(par_done_reg693_done)
  );
  
  std_reg #(1) par_done_reg694 (
      .in(par_done_reg694_in),
      .write_en(par_done_reg694_write_en),
      .clk(clk),
      .out(par_done_reg694_out),
      .done(par_done_reg694_done)
  );
  
  std_reg #(1) par_done_reg695 (
      .in(par_done_reg695_in),
      .write_en(par_done_reg695_write_en),
      .clk(clk),
      .out(par_done_reg695_out),
      .done(par_done_reg695_done)
  );
  
  std_reg #(1) par_done_reg696 (
      .in(par_done_reg696_in),
      .write_en(par_done_reg696_write_en),
      .clk(clk),
      .out(par_done_reg696_out),
      .done(par_done_reg696_done)
  );
  
  std_reg #(1) par_done_reg697 (
      .in(par_done_reg697_in),
      .write_en(par_done_reg697_write_en),
      .clk(clk),
      .out(par_done_reg697_out),
      .done(par_done_reg697_done)
  );
  
  std_reg #(1) par_done_reg698 (
      .in(par_done_reg698_in),
      .write_en(par_done_reg698_write_en),
      .clk(clk),
      .out(par_done_reg698_out),
      .done(par_done_reg698_done)
  );
  
  std_reg #(1) par_done_reg699 (
      .in(par_done_reg699_in),
      .write_en(par_done_reg699_write_en),
      .clk(clk),
      .out(par_done_reg699_out),
      .done(par_done_reg699_done)
  );
  
  std_reg #(1) par_done_reg700 (
      .in(par_done_reg700_in),
      .write_en(par_done_reg700_write_en),
      .clk(clk),
      .out(par_done_reg700_out),
      .done(par_done_reg700_done)
  );
  
  std_reg #(1) par_done_reg701 (
      .in(par_done_reg701_in),
      .write_en(par_done_reg701_write_en),
      .clk(clk),
      .out(par_done_reg701_out),
      .done(par_done_reg701_done)
  );
  
  std_reg #(1) par_reset28 (
      .in(par_reset28_in),
      .write_en(par_reset28_write_en),
      .clk(clk),
      .out(par_reset28_out),
      .done(par_reset28_done)
  );
  
  std_reg #(1) par_done_reg702 (
      .in(par_done_reg702_in),
      .write_en(par_done_reg702_write_en),
      .clk(clk),
      .out(par_done_reg702_out),
      .done(par_done_reg702_done)
  );
  
  std_reg #(1) par_done_reg703 (
      .in(par_done_reg703_in),
      .write_en(par_done_reg703_write_en),
      .clk(clk),
      .out(par_done_reg703_out),
      .done(par_done_reg703_done)
  );
  
  std_reg #(1) par_done_reg704 (
      .in(par_done_reg704_in),
      .write_en(par_done_reg704_write_en),
      .clk(clk),
      .out(par_done_reg704_out),
      .done(par_done_reg704_done)
  );
  
  std_reg #(1) par_done_reg705 (
      .in(par_done_reg705_in),
      .write_en(par_done_reg705_write_en),
      .clk(clk),
      .out(par_done_reg705_out),
      .done(par_done_reg705_done)
  );
  
  std_reg #(1) par_done_reg706 (
      .in(par_done_reg706_in),
      .write_en(par_done_reg706_write_en),
      .clk(clk),
      .out(par_done_reg706_out),
      .done(par_done_reg706_done)
  );
  
  std_reg #(1) par_done_reg707 (
      .in(par_done_reg707_in),
      .write_en(par_done_reg707_write_en),
      .clk(clk),
      .out(par_done_reg707_out),
      .done(par_done_reg707_done)
  );
  
  std_reg #(1) par_done_reg708 (
      .in(par_done_reg708_in),
      .write_en(par_done_reg708_write_en),
      .clk(clk),
      .out(par_done_reg708_out),
      .done(par_done_reg708_done)
  );
  
  std_reg #(1) par_done_reg709 (
      .in(par_done_reg709_in),
      .write_en(par_done_reg709_write_en),
      .clk(clk),
      .out(par_done_reg709_out),
      .done(par_done_reg709_done)
  );
  
  std_reg #(1) par_done_reg710 (
      .in(par_done_reg710_in),
      .write_en(par_done_reg710_write_en),
      .clk(clk),
      .out(par_done_reg710_out),
      .done(par_done_reg710_done)
  );
  
  std_reg #(1) par_done_reg711 (
      .in(par_done_reg711_in),
      .write_en(par_done_reg711_write_en),
      .clk(clk),
      .out(par_done_reg711_out),
      .done(par_done_reg711_done)
  );
  
  std_reg #(1) par_done_reg712 (
      .in(par_done_reg712_in),
      .write_en(par_done_reg712_write_en),
      .clk(clk),
      .out(par_done_reg712_out),
      .done(par_done_reg712_done)
  );
  
  std_reg #(1) par_done_reg713 (
      .in(par_done_reg713_in),
      .write_en(par_done_reg713_write_en),
      .clk(clk),
      .out(par_done_reg713_out),
      .done(par_done_reg713_done)
  );
  
  std_reg #(1) par_reset29 (
      .in(par_reset29_in),
      .write_en(par_reset29_write_en),
      .clk(clk),
      .out(par_reset29_out),
      .done(par_reset29_done)
  );
  
  std_reg #(1) par_done_reg714 (
      .in(par_done_reg714_in),
      .write_en(par_done_reg714_write_en),
      .clk(clk),
      .out(par_done_reg714_out),
      .done(par_done_reg714_done)
  );
  
  std_reg #(1) par_done_reg715 (
      .in(par_done_reg715_in),
      .write_en(par_done_reg715_write_en),
      .clk(clk),
      .out(par_done_reg715_out),
      .done(par_done_reg715_done)
  );
  
  std_reg #(1) par_done_reg716 (
      .in(par_done_reg716_in),
      .write_en(par_done_reg716_write_en),
      .clk(clk),
      .out(par_done_reg716_out),
      .done(par_done_reg716_done)
  );
  
  std_reg #(1) par_done_reg717 (
      .in(par_done_reg717_in),
      .write_en(par_done_reg717_write_en),
      .clk(clk),
      .out(par_done_reg717_out),
      .done(par_done_reg717_done)
  );
  
  std_reg #(1) par_done_reg718 (
      .in(par_done_reg718_in),
      .write_en(par_done_reg718_write_en),
      .clk(clk),
      .out(par_done_reg718_out),
      .done(par_done_reg718_done)
  );
  
  std_reg #(1) par_done_reg719 (
      .in(par_done_reg719_in),
      .write_en(par_done_reg719_write_en),
      .clk(clk),
      .out(par_done_reg719_out),
      .done(par_done_reg719_done)
  );
  
  std_reg #(1) par_reset30 (
      .in(par_reset30_in),
      .write_en(par_reset30_write_en),
      .clk(clk),
      .out(par_reset30_out),
      .done(par_reset30_done)
  );
  
  std_reg #(1) par_done_reg720 (
      .in(par_done_reg720_in),
      .write_en(par_done_reg720_write_en),
      .clk(clk),
      .out(par_done_reg720_out),
      .done(par_done_reg720_done)
  );
  
  std_reg #(1) par_done_reg721 (
      .in(par_done_reg721_in),
      .write_en(par_done_reg721_write_en),
      .clk(clk),
      .out(par_done_reg721_out),
      .done(par_done_reg721_done)
  );
  
  std_reg #(1) par_done_reg722 (
      .in(par_done_reg722_in),
      .write_en(par_done_reg722_write_en),
      .clk(clk),
      .out(par_done_reg722_out),
      .done(par_done_reg722_done)
  );
  
  std_reg #(1) par_done_reg723 (
      .in(par_done_reg723_in),
      .write_en(par_done_reg723_write_en),
      .clk(clk),
      .out(par_done_reg723_out),
      .done(par_done_reg723_done)
  );
  
  std_reg #(1) par_done_reg724 (
      .in(par_done_reg724_in),
      .write_en(par_done_reg724_write_en),
      .clk(clk),
      .out(par_done_reg724_out),
      .done(par_done_reg724_done)
  );
  
  std_reg #(1) par_done_reg725 (
      .in(par_done_reg725_in),
      .write_en(par_done_reg725_write_en),
      .clk(clk),
      .out(par_done_reg725_out),
      .done(par_done_reg725_done)
  );
  
  std_reg #(1) par_reset31 (
      .in(par_reset31_in),
      .write_en(par_reset31_write_en),
      .clk(clk),
      .out(par_reset31_out),
      .done(par_reset31_done)
  );
  
  std_reg #(1) par_done_reg726 (
      .in(par_done_reg726_in),
      .write_en(par_done_reg726_write_en),
      .clk(clk),
      .out(par_done_reg726_out),
      .done(par_done_reg726_done)
  );
  
  std_reg #(1) par_done_reg727 (
      .in(par_done_reg727_in),
      .write_en(par_done_reg727_write_en),
      .clk(clk),
      .out(par_done_reg727_out),
      .done(par_done_reg727_done)
  );
  
  std_reg #(1) par_done_reg728 (
      .in(par_done_reg728_in),
      .write_en(par_done_reg728_write_en),
      .clk(clk),
      .out(par_done_reg728_out),
      .done(par_done_reg728_done)
  );
  
  std_reg #(1) par_reset32 (
      .in(par_reset32_in),
      .write_en(par_reset32_write_en),
      .clk(clk),
      .out(par_reset32_out),
      .done(par_reset32_done)
  );
  
  std_reg #(1) par_done_reg729 (
      .in(par_done_reg729_in),
      .write_en(par_done_reg729_write_en),
      .clk(clk),
      .out(par_done_reg729_out),
      .done(par_done_reg729_done)
  );
  
  std_reg #(1) par_done_reg730 (
      .in(par_done_reg730_in),
      .write_en(par_done_reg730_write_en),
      .clk(clk),
      .out(par_done_reg730_out),
      .done(par_done_reg730_done)
  );
  
  std_reg #(1) par_reset33 (
      .in(par_reset33_in),
      .write_en(par_reset33_write_en),
      .clk(clk),
      .out(par_reset33_out),
      .done(par_reset33_done)
  );
  
  std_reg #(1) par_done_reg731 (
      .in(par_done_reg731_in),
      .write_en(par_done_reg731_write_en),
      .clk(clk),
      .out(par_done_reg731_out),
      .done(par_done_reg731_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign done = (fsm0_out == 32'd70) ? 1'd1 : '0;
  assign out_mem_addr0 = (fsm0_out == 32'd64 & !out_mem_done & go | fsm0_out == 32'd65 & !out_mem_done & go | fsm0_out == 32'd66 & !out_mem_done & go | fsm0_out == 32'd67 & !out_mem_done & go | fsm0_out == 32'd68 & !out_mem_done & go | fsm0_out == 32'd69 & !out_mem_done & go) ? 3'd5 : (fsm0_out == 32'd58 & !out_mem_done & go | fsm0_out == 32'd59 & !out_mem_done & go | fsm0_out == 32'd60 & !out_mem_done & go | fsm0_out == 32'd61 & !out_mem_done & go | fsm0_out == 32'd62 & !out_mem_done & go | fsm0_out == 32'd63 & !out_mem_done & go) ? 3'd4 : (fsm0_out == 32'd52 & !out_mem_done & go | fsm0_out == 32'd53 & !out_mem_done & go | fsm0_out == 32'd54 & !out_mem_done & go | fsm0_out == 32'd55 & !out_mem_done & go | fsm0_out == 32'd56 & !out_mem_done & go | fsm0_out == 32'd57 & !out_mem_done & go) ? 3'd3 : (fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go) ? 3'd2 : (fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go | fsm0_out == 32'd38 & !out_mem_done & go | fsm0_out == 32'd39 & !out_mem_done & go) ? 3'd0 : (fsm0_out == 32'd40 & !out_mem_done & go | fsm0_out == 32'd41 & !out_mem_done & go | fsm0_out == 32'd42 & !out_mem_done & go | fsm0_out == 32'd43 & !out_mem_done & go | fsm0_out == 32'd44 & !out_mem_done & go | fsm0_out == 32'd45 & !out_mem_done & go) ? 3'd1 : '0;
  assign out_mem_addr1 = (fsm0_out == 32'd39 & !out_mem_done & go | fsm0_out == 32'd45 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd57 & !out_mem_done & go | fsm0_out == 32'd63 & !out_mem_done & go | fsm0_out == 32'd69 & !out_mem_done & go) ? 3'd5 : (fsm0_out == 32'd38 & !out_mem_done & go | fsm0_out == 32'd44 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd56 & !out_mem_done & go | fsm0_out == 32'd62 & !out_mem_done & go | fsm0_out == 32'd68 & !out_mem_done & go) ? 3'd4 : (fsm0_out == 32'd37 & !out_mem_done & go | fsm0_out == 32'd43 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd55 & !out_mem_done & go | fsm0_out == 32'd61 & !out_mem_done & go | fsm0_out == 32'd67 & !out_mem_done & go) ? 3'd3 : (fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd42 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd54 & !out_mem_done & go | fsm0_out == 32'd60 & !out_mem_done & go | fsm0_out == 32'd66 & !out_mem_done & go) ? 3'd2 : (fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd40 & !out_mem_done & go | fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go | fsm0_out == 32'd58 & !out_mem_done & go | fsm0_out == 32'd64 & !out_mem_done & go) ? 3'd0 : (fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd41 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd53 & !out_mem_done & go | fsm0_out == 32'd59 & !out_mem_done & go | fsm0_out == 32'd65 & !out_mem_done & go) ? 3'd1 : '0;
  assign out_mem_write_data = (fsm0_out == 32'd69 & !out_mem_done & go) ? pe_55_out : (fsm0_out == 32'd68 & !out_mem_done & go) ? pe_54_out : (fsm0_out == 32'd67 & !out_mem_done & go) ? pe_53_out : (fsm0_out == 32'd66 & !out_mem_done & go) ? pe_52_out : (fsm0_out == 32'd65 & !out_mem_done & go) ? pe_51_out : (fsm0_out == 32'd64 & !out_mem_done & go) ? pe_50_out : (fsm0_out == 32'd63 & !out_mem_done & go) ? pe_45_out : (fsm0_out == 32'd62 & !out_mem_done & go) ? pe_44_out : (fsm0_out == 32'd61 & !out_mem_done & go) ? pe_43_out : (fsm0_out == 32'd60 & !out_mem_done & go) ? pe_42_out : (fsm0_out == 32'd59 & !out_mem_done & go) ? pe_41_out : (fsm0_out == 32'd58 & !out_mem_done & go) ? pe_40_out : (fsm0_out == 32'd57 & !out_mem_done & go) ? pe_35_out : (fsm0_out == 32'd56 & !out_mem_done & go) ? pe_34_out : (fsm0_out == 32'd55 & !out_mem_done & go) ? pe_33_out : (fsm0_out == 32'd54 & !out_mem_done & go) ? pe_32_out : (fsm0_out == 32'd53 & !out_mem_done & go) ? pe_31_out : (fsm0_out == 32'd52 & !out_mem_done & go) ? pe_30_out : (fsm0_out == 32'd51 & !out_mem_done & go) ? pe_25_out : (fsm0_out == 32'd50 & !out_mem_done & go) ? pe_24_out : (fsm0_out == 32'd49 & !out_mem_done & go) ? pe_23_out : (fsm0_out == 32'd48 & !out_mem_done & go) ? pe_22_out : (fsm0_out == 32'd47 & !out_mem_done & go) ? pe_21_out : (fsm0_out == 32'd46 & !out_mem_done & go) ? pe_20_out : (fsm0_out == 32'd45 & !out_mem_done & go) ? pe_15_out : (fsm0_out == 32'd44 & !out_mem_done & go) ? pe_14_out : (fsm0_out == 32'd43 & !out_mem_done & go) ? pe_13_out : (fsm0_out == 32'd42 & !out_mem_done & go) ? pe_12_out : (fsm0_out == 32'd41 & !out_mem_done & go) ? pe_11_out : (fsm0_out == 32'd40 & !out_mem_done & go) ? pe_10_out : (fsm0_out == 32'd39 & !out_mem_done & go) ? pe_05_out : (fsm0_out == 32'd38 & !out_mem_done & go) ? pe_04_out : (fsm0_out == 32'd37 & !out_mem_done & go) ? pe_03_out : (fsm0_out == 32'd36 & !out_mem_done & go) ? pe_02_out : (fsm0_out == 32'd35 & !out_mem_done & go) ? pe_01_out : (fsm0_out == 32'd34 & !out_mem_done & go) ? pe_00_out : '0;
  assign out_mem_write_en = (fsm0_out == 32'd34 & !out_mem_done & go | fsm0_out == 32'd35 & !out_mem_done & go | fsm0_out == 32'd36 & !out_mem_done & go | fsm0_out == 32'd37 & !out_mem_done & go | fsm0_out == 32'd38 & !out_mem_done & go | fsm0_out == 32'd39 & !out_mem_done & go | fsm0_out == 32'd40 & !out_mem_done & go | fsm0_out == 32'd41 & !out_mem_done & go | fsm0_out == 32'd42 & !out_mem_done & go | fsm0_out == 32'd43 & !out_mem_done & go | fsm0_out == 32'd44 & !out_mem_done & go | fsm0_out == 32'd45 & !out_mem_done & go | fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go | fsm0_out == 32'd53 & !out_mem_done & go | fsm0_out == 32'd54 & !out_mem_done & go | fsm0_out == 32'd55 & !out_mem_done & go | fsm0_out == 32'd56 & !out_mem_done & go | fsm0_out == 32'd57 & !out_mem_done & go | fsm0_out == 32'd58 & !out_mem_done & go | fsm0_out == 32'd59 & !out_mem_done & go | fsm0_out == 32'd60 & !out_mem_done & go | fsm0_out == 32'd61 & !out_mem_done & go | fsm0_out == 32'd62 & !out_mem_done & go | fsm0_out == 32'd63 & !out_mem_done & go | fsm0_out == 32'd64 & !out_mem_done & go | fsm0_out == 32'd65 & !out_mem_done & go | fsm0_out == 32'd66 & !out_mem_done & go | fsm0_out == 32'd67 & !out_mem_done & go | fsm0_out == 32'd68 & !out_mem_done & go | fsm0_out == 32'd69 & !out_mem_done & go) ? 1'd1 : '0;
  assign left_55_read_in = (!(par_done_reg605_out | left_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg656_out | left_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg691_out | left_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg713_out | left_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg725_out | left_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg730_out | left_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_54_write_out : '0;
  assign left_55_read_write_en = (!(par_done_reg605_out | left_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg656_out | left_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg691_out | left_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg713_out | left_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg725_out | left_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg730_out | left_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_55_read_in = (!(par_done_reg584_out | top_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg641_out | top_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg681_out | top_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg707_out | top_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg722_out | top_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg729_out | top_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_45_write_out : '0;
  assign top_55_read_write_en = (!(par_done_reg584_out | top_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg641_out | top_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg681_out | top_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg707_out | top_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg722_out | top_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg729_out | top_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_55_top = (!(par_done_reg626_out | pe_55_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg671_out | pe_55_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg701_out | pe_55_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg719_out | pe_55_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg728_out | pe_55_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg731_out | pe_55_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_55_read_out : '0;
  assign pe_55_left = (!(par_done_reg626_out | pe_55_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg671_out | pe_55_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg701_out | pe_55_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg719_out | pe_55_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg728_out | pe_55_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg731_out | pe_55_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_55_read_out : '0;
  assign pe_55_go = (!pe_55_done & (!(par_done_reg626_out | pe_55_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg671_out | pe_55_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg701_out | pe_55_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg719_out | pe_55_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg728_out | pe_55_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg731_out | pe_55_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_54_write_in = (pe_54_done & (!(par_done_reg563_out | right_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg625_out | right_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg670_out | right_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg700_out | right_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg718_out | right_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg727_out | right_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_54_right : '0;
  assign right_54_write_write_en = (pe_54_done & (!(par_done_reg563_out | right_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg625_out | right_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg670_out | right_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg700_out | right_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg718_out | right_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg727_out | right_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_54_read_in = (!(par_done_reg536_out | left_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg604_out | left_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg655_out | left_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg690_out | left_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg712_out | left_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg724_out | left_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_53_write_out : '0;
  assign left_54_read_write_en = (!(par_done_reg536_out | left_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg604_out | left_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg655_out | left_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg690_out | left_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg712_out | left_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg724_out | left_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_54_read_in = (!(par_done_reg511_out | top_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg583_out | top_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg640_out | top_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg680_out | top_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg706_out | top_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg721_out | top_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_44_write_out : '0;
  assign top_54_read_write_en = (!(par_done_reg511_out | top_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg583_out | top_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg640_out | top_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg680_out | top_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg706_out | top_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg721_out | top_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_54_top = (!(par_done_reg563_out | right_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg625_out | right_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg670_out | right_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg700_out | right_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg718_out | right_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg727_out | right_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_54_read_out : '0;
  assign pe_54_left = (!(par_done_reg563_out | right_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg625_out | right_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg670_out | right_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg700_out | right_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg718_out | right_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg727_out | right_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_54_read_out : '0;
  assign pe_54_go = (!pe_54_done & (!(par_done_reg563_out | right_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg625_out | right_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg670_out | right_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg700_out | right_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg718_out | right_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg727_out | right_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_53_write_in = (pe_53_done & (!(par_done_reg486_out | right_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg562_out | right_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg624_out | right_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg669_out | right_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg699_out | right_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg717_out | right_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_53_right : '0;
  assign right_53_write_write_en = (pe_53_done & (!(par_done_reg486_out | right_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg562_out | right_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg624_out | right_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg669_out | right_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg699_out | right_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg717_out | right_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_53_read_in = (!(par_done_reg455_out | left_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg535_out | left_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg603_out | left_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg654_out | left_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg689_out | left_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg711_out | left_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_52_write_out : '0;
  assign left_53_read_write_en = (!(par_done_reg455_out | left_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg535_out | left_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg603_out | left_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg654_out | left_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg689_out | left_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg711_out | left_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_53_read_in = (!(par_done_reg428_out | top_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg510_out | top_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg582_out | top_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg639_out | top_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg679_out | top_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg705_out | top_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_43_write_out : '0;
  assign top_53_read_write_en = (!(par_done_reg428_out | top_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg510_out | top_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg582_out | top_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg639_out | top_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg679_out | top_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg705_out | top_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_53_top = (!(par_done_reg486_out | right_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg562_out | right_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg624_out | right_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg669_out | right_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg699_out | right_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg717_out | right_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_53_read_out : '0;
  assign pe_53_left = (!(par_done_reg486_out | right_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg562_out | right_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg624_out | right_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg669_out | right_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg699_out | right_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg717_out | right_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_53_read_out : '0;
  assign pe_53_go = (!pe_53_done & (!(par_done_reg486_out | right_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg562_out | right_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg624_out | right_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg669_out | right_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg699_out | right_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg717_out | right_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_52_write_in = (pe_52_done & (!(par_done_reg401_out | right_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg485_out | right_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg561_out | right_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg623_out | right_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg668_out | right_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg698_out | right_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_52_right : '0;
  assign right_52_write_write_en = (pe_52_done & (!(par_done_reg401_out | right_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg485_out | right_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg561_out | right_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg623_out | right_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg668_out | right_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg698_out | right_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_52_read_in = (!(par_done_reg368_out | left_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg454_out | left_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg534_out | left_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg602_out | left_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg653_out | left_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg688_out | left_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_51_write_out : '0;
  assign left_52_read_write_en = (!(par_done_reg368_out | left_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg454_out | left_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg534_out | left_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg602_out | left_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg653_out | left_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg688_out | left_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_52_read_in = (!(par_done_reg341_out | top_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg427_out | top_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg509_out | top_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg581_out | top_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg638_out | top_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg678_out | top_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_42_write_out : '0;
  assign top_52_read_write_en = (!(par_done_reg341_out | top_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg427_out | top_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg509_out | top_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg581_out | top_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg638_out | top_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg678_out | top_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_52_top = (!(par_done_reg401_out | right_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg485_out | right_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg561_out | right_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg623_out | right_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg668_out | right_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg698_out | right_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_52_read_out : '0;
  assign pe_52_left = (!(par_done_reg401_out | right_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg485_out | right_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg561_out | right_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg623_out | right_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg668_out | right_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg698_out | right_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_52_read_out : '0;
  assign pe_52_go = (!pe_52_done & (!(par_done_reg401_out | right_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg485_out | right_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg561_out | right_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg623_out | right_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg668_out | right_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg698_out | right_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_51_write_in = (pe_51_done & (!(par_done_reg314_out | right_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg400_out | right_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg484_out | right_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg560_out | right_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg622_out | right_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg667_out | right_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_51_right : '0;
  assign right_51_write_write_en = (pe_51_done & (!(par_done_reg314_out | right_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg400_out | right_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg484_out | right_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg560_out | right_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg622_out | right_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg667_out | right_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_51_read_in = (!(par_done_reg281_out | left_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg367_out | left_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg453_out | left_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg533_out | left_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg601_out | left_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg652_out | left_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_50_write_out : '0;
  assign left_51_read_write_en = (!(par_done_reg281_out | left_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg367_out | left_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg453_out | left_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg533_out | left_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg601_out | left_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg652_out | left_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_51_read_in = (!(par_done_reg256_out | top_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg340_out | top_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg426_out | top_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg508_out | top_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg580_out | top_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg637_out | top_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_41_write_out : '0;
  assign top_51_read_write_en = (!(par_done_reg256_out | top_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg340_out | top_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg426_out | top_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg508_out | top_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg580_out | top_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg637_out | top_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_51_top = (!(par_done_reg314_out | right_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg400_out | right_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg484_out | right_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg560_out | right_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg622_out | right_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg667_out | right_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_51_read_out : '0;
  assign pe_51_left = (!(par_done_reg314_out | right_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg400_out | right_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg484_out | right_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg560_out | right_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg622_out | right_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg667_out | right_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_51_read_out : '0;
  assign pe_51_go = (!pe_51_done & (!(par_done_reg314_out | right_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg400_out | right_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg484_out | right_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg560_out | right_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg622_out | right_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg667_out | right_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_50_write_in = (pe_50_done & (!(par_done_reg231_out | right_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg399_out | right_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg483_out | right_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg559_out | right_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg621_out | right_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_50_right : '0;
  assign right_50_write_write_en = (pe_50_done & (!(par_done_reg231_out | right_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg399_out | right_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg483_out | right_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg559_out | right_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg621_out | right_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_50_read_in = (!(par_done_reg200_out | left_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg280_out | left_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg366_out | left_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg452_out | left_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg532_out | left_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg600_out | left_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? l5_read_data : '0;
  assign left_50_read_write_en = (!(par_done_reg200_out | left_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg280_out | left_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg366_out | left_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg452_out | left_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg532_out | left_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg600_out | left_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_50_read_in = (!(par_done_reg179_out | top_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg255_out | top_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg339_out | top_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg425_out | top_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg507_out | top_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg579_out | top_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_40_write_out : '0;
  assign top_50_read_write_en = (!(par_done_reg179_out | top_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg255_out | top_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg339_out | top_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg425_out | top_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg507_out | top_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg579_out | top_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_50_top = (!(par_done_reg231_out | right_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg399_out | right_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg483_out | right_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg559_out | right_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg621_out | right_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_50_read_out : '0;
  assign pe_50_left = (!(par_done_reg231_out | right_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg399_out | right_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg483_out | right_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg559_out | right_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg621_out | right_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_50_read_out : '0;
  assign pe_50_go = (!pe_50_done & (!(par_done_reg231_out | right_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg399_out | right_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg483_out | right_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg559_out | right_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg621_out | right_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_45_write_in = (pe_45_done & (!(par_done_reg558_out | down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg620_out | down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg666_out | down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg697_out | down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg716_out | down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg726_out | down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_45_down : '0;
  assign down_45_write_write_en = (pe_45_done & (!(par_done_reg558_out | down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg620_out | down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg666_out | down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg697_out | down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg716_out | down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg726_out | down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_45_read_in = (!(par_done_reg531_out | left_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg599_out | left_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg651_out | left_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg687_out | left_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg710_out | left_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg723_out | left_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_44_write_out : '0;
  assign left_45_read_write_en = (!(par_done_reg531_out | left_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg599_out | left_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg651_out | left_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg687_out | left_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg710_out | left_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg723_out | left_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_45_read_in = (!(par_done_reg506_out | top_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg578_out | top_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg636_out | top_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg677_out | top_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg704_out | top_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg720_out | top_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_35_write_out : '0;
  assign top_45_read_write_en = (!(par_done_reg506_out | top_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg578_out | top_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg636_out | top_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg677_out | top_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg704_out | top_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg720_out | top_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_45_top = (!(par_done_reg558_out | down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg620_out | down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg666_out | down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg697_out | down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg716_out | down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg726_out | down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_45_read_out : '0;
  assign pe_45_left = (!(par_done_reg558_out | down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg620_out | down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg666_out | down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg697_out | down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg716_out | down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg726_out | down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_45_read_out : '0;
  assign pe_45_go = (!pe_45_done & (!(par_done_reg558_out | down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg620_out | down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg666_out | down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg697_out | down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg716_out | down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg726_out | down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_44_write_in = (pe_44_done & (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_44_down : '0;
  assign down_44_write_write_en = (pe_44_done & (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_44_write_in = (pe_44_done & (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_44_right : '0;
  assign right_44_write_write_en = (pe_44_done & (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_44_read_in = (!(par_done_reg451_out | left_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg530_out | left_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg598_out | left_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg650_out | left_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg686_out | left_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg709_out | left_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_43_write_out : '0;
  assign left_44_read_write_en = (!(par_done_reg451_out | left_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg530_out | left_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg598_out | left_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg650_out | left_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg686_out | left_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg709_out | left_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_44_read_in = (!(par_done_reg424_out | top_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg505_out | top_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg577_out | top_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg635_out | top_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg676_out | top_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg703_out | top_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_34_write_out : '0;
  assign top_44_read_write_en = (!(par_done_reg424_out | top_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg505_out | top_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg577_out | top_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg635_out | top_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg676_out | top_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg703_out | top_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_44_top = (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_44_read_out : '0;
  assign pe_44_left = (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_44_read_out : '0;
  assign pe_44_go = (!pe_44_done & (!(par_done_reg482_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg557_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg619_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg665_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg696_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg715_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_43_write_in = (pe_43_done & (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_43_down : '0;
  assign down_43_write_write_en = (pe_43_done & (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_43_write_in = (pe_43_done & (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_43_right : '0;
  assign right_43_write_write_en = (pe_43_done & (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_43_read_in = (!(par_done_reg365_out | left_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg450_out | left_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg529_out | left_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg597_out | left_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg649_out | left_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg685_out | left_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_42_write_out : '0;
  assign left_43_read_write_en = (!(par_done_reg365_out | left_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg450_out | left_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg529_out | left_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg597_out | left_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg649_out | left_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg685_out | left_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_43_read_in = (!(par_done_reg338_out | top_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg423_out | top_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg504_out | top_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg576_out | top_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg634_out | top_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg675_out | top_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_33_write_out : '0;
  assign top_43_read_write_en = (!(par_done_reg338_out | top_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg423_out | top_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg504_out | top_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg576_out | top_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg634_out | top_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg675_out | top_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_43_top = (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_43_read_out : '0;
  assign pe_43_left = (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_43_read_out : '0;
  assign pe_43_go = (!pe_43_done & (!(par_done_reg398_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg481_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg556_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg618_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg664_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg695_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_42_write_in = (pe_42_done & (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_42_down : '0;
  assign down_42_write_write_en = (pe_42_done & (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_42_write_in = (pe_42_done & (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_42_right : '0;
  assign right_42_write_write_en = (pe_42_done & (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_42_read_in = (!(par_done_reg279_out | left_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg364_out | left_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg449_out | left_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg528_out | left_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg596_out | left_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg648_out | left_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_41_write_out : '0;
  assign left_42_read_write_en = (!(par_done_reg279_out | left_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg364_out | left_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg449_out | left_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg528_out | left_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg596_out | left_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg648_out | left_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_42_read_in = (!(par_done_reg254_out | top_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg337_out | top_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg422_out | top_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg503_out | top_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg575_out | top_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg633_out | top_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_32_write_out : '0;
  assign top_42_read_write_en = (!(par_done_reg254_out | top_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg337_out | top_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg422_out | top_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg503_out | top_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg575_out | top_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg633_out | top_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_42_top = (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_42_read_out : '0;
  assign pe_42_left = (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_42_read_out : '0;
  assign pe_42_go = (!pe_42_done & (!(par_done_reg312_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg397_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg480_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg555_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg617_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg663_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_41_write_in = (pe_41_done & (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_41_down : '0;
  assign down_41_write_write_en = (pe_41_done & (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_41_write_in = (pe_41_done & (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_41_right : '0;
  assign right_41_write_write_en = (pe_41_done & (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_41_read_in = (!(par_done_reg199_out | left_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg278_out | left_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg363_out | left_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg448_out | left_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg527_out | left_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg595_out | left_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_40_write_out : '0;
  assign left_41_read_write_en = (!(par_done_reg199_out | left_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg278_out | left_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg363_out | left_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg448_out | left_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg527_out | left_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg595_out | left_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_41_read_in = (!(par_done_reg178_out | top_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg253_out | top_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg336_out | top_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg421_out | top_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg502_out | top_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg574_out | top_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_31_write_out : '0;
  assign top_41_read_write_en = (!(par_done_reg178_out | top_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg253_out | top_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg336_out | top_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg421_out | top_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg502_out | top_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg574_out | top_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_41_top = (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_41_read_out : '0;
  assign pe_41_left = (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_41_read_out : '0;
  assign pe_41_go = (!pe_41_done & (!(par_done_reg230_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg311_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg396_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg479_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg554_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg616_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_40_write_in = (pe_40_done & (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_40_down : '0;
  assign down_40_write_write_en = (pe_40_done & (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_40_write_in = (pe_40_done & (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_40_right : '0;
  assign right_40_write_write_en = (pe_40_done & (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_40_read_in = (!(par_done_reg131_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg198_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg277_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg362_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg447_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg526_out | left_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? l4_read_data : '0;
  assign left_40_read_write_en = (!(par_done_reg131_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg198_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg277_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg362_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg447_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg526_out | left_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_40_read_in = (!(par_done_reg116_out | top_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg177_out | top_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg252_out | top_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg335_out | top_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg420_out | top_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg501_out | top_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_30_write_out : '0;
  assign top_40_read_write_en = (!(par_done_reg116_out | top_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg177_out | top_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg252_out | top_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg335_out | top_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg420_out | top_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg501_out | top_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_40_top = (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_40_read_out : '0;
  assign pe_40_left = (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_40_read_out : '0;
  assign pe_40_go = (!pe_40_done & (!(par_done_reg158_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg229_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg395_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg478_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg553_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_35_write_in = (pe_35_done & (!(par_done_reg477_out | down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg552_out | down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg615_out | down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg662_out | down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg694_out | down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg714_out | down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_35_down : '0;
  assign down_35_write_write_en = (pe_35_done & (!(par_done_reg477_out | down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg552_out | down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg615_out | down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg662_out | down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg694_out | down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg714_out | down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_35_read_in = (!(par_done_reg446_out | left_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg525_out | left_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg594_out | left_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg647_out | left_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg684_out | left_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg708_out | left_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_34_write_out : '0;
  assign left_35_read_write_en = (!(par_done_reg446_out | left_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg525_out | left_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg594_out | left_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg647_out | left_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg684_out | left_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg708_out | left_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_35_read_in = (!(par_done_reg419_out | top_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg500_out | top_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg573_out | top_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg632_out | top_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg674_out | top_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg702_out | top_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_25_write_out : '0;
  assign top_35_read_write_en = (!(par_done_reg419_out | top_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg500_out | top_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg573_out | top_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg632_out | top_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg674_out | top_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg702_out | top_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_35_top = (!(par_done_reg477_out | down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg552_out | down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg615_out | down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg662_out | down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg694_out | down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg714_out | down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_35_read_out : '0;
  assign pe_35_left = (!(par_done_reg477_out | down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg552_out | down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg615_out | down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg662_out | down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg694_out | down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg714_out | down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_35_read_out : '0;
  assign pe_35_go = (!pe_35_done & (!(par_done_reg477_out | down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg552_out | down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg615_out | down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg662_out | down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg694_out | down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg714_out | down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_34_write_in = (pe_34_done & (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_34_down : '0;
  assign down_34_write_write_en = (pe_34_done & (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_34_write_in = (pe_34_done & (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_34_right : '0;
  assign right_34_write_write_en = (pe_34_done & (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_34_read_in = (!(par_done_reg361_out | left_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg445_out | left_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg524_out | left_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg593_out | left_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg646_out | left_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg683_out | left_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_33_write_out : '0;
  assign left_34_read_write_en = (!(par_done_reg361_out | left_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg445_out | left_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg524_out | left_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg593_out | left_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg646_out | left_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg683_out | left_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_34_read_in = (!(par_done_reg334_out | top_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg418_out | top_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg499_out | top_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg572_out | top_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg631_out | top_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg673_out | top_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_24_write_out : '0;
  assign top_34_read_write_en = (!(par_done_reg334_out | top_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg418_out | top_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg499_out | top_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg572_out | top_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg631_out | top_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg673_out | top_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_34_top = (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_34_read_out : '0;
  assign pe_34_left = (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_34_read_out : '0;
  assign pe_34_go = (!pe_34_done & (!(par_done_reg394_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg476_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg551_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg614_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg661_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg693_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_33_write_in = (pe_33_done & (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_33_down : '0;
  assign down_33_write_write_en = (pe_33_done & (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_33_write_in = (pe_33_done & (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_33_right : '0;
  assign right_33_write_write_en = (pe_33_done & (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_33_read_in = (!(par_done_reg276_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg360_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg444_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg523_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg592_out | left_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg645_out | left_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_32_write_out : '0;
  assign left_33_read_write_en = (!(par_done_reg276_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg360_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg444_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg523_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg592_out | left_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg645_out | left_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_33_read_in = (!(par_done_reg251_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg333_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg417_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg498_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg571_out | top_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg630_out | top_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_23_write_out : '0;
  assign top_33_read_write_en = (!(par_done_reg251_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg333_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg417_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg498_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg571_out | top_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg630_out | top_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_33_top = (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_33_read_out : '0;
  assign pe_33_left = (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_33_read_out : '0;
  assign pe_33_go = (!pe_33_done & (!(par_done_reg309_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg393_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg475_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg550_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg613_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg660_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_32_write_in = (pe_32_done & (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_32_down : '0;
  assign down_32_write_write_en = (pe_32_done & (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_32_write_in = (pe_32_done & (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_32_right : '0;
  assign right_32_write_write_en = (pe_32_done & (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_32_read_in = (!(par_done_reg197_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg275_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg359_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg443_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg522_out | left_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg591_out | left_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_31_write_out : '0;
  assign left_32_read_write_en = (!(par_done_reg197_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg275_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg359_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg443_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg522_out | left_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg591_out | left_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_32_read_in = (!(par_done_reg176_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg250_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg332_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg416_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg497_out | top_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg570_out | top_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_22_write_out : '0;
  assign top_32_read_write_en = (!(par_done_reg176_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg250_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg332_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg416_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg497_out | top_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg570_out | top_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_32_top = (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_32_read_out : '0;
  assign pe_32_left = (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_32_read_out : '0;
  assign pe_32_go = (!pe_32_done & (!(par_done_reg228_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg392_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg474_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg549_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg612_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_31_write_in = (pe_31_done & (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_31_down : '0;
  assign down_31_write_write_en = (pe_31_done & (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_31_write_in = (pe_31_done & (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_31_right : '0;
  assign right_31_write_write_en = (pe_31_done & (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_31_read_in = (!(par_done_reg130_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg196_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg274_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg358_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg442_out | left_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg521_out | left_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_30_write_out : '0;
  assign left_31_read_write_en = (!(par_done_reg130_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg196_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg274_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg358_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg442_out | left_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg521_out | left_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_31_read_in = (!(par_done_reg115_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg249_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg331_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg415_out | top_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg496_out | top_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_21_write_out : '0;
  assign top_31_read_write_en = (!(par_done_reg115_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg249_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg331_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg415_out | top_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg496_out | top_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_31_top = (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_31_read_out : '0;
  assign pe_31_left = (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_31_read_out : '0;
  assign pe_31_go = (!pe_31_done & (!(par_done_reg157_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg391_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg473_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg548_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_30_write_in = (pe_30_done & (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_30_down : '0;
  assign down_30_write_write_en = (pe_30_done & (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_30_write_in = (pe_30_done & (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_30_right : '0;
  assign right_30_write_write_en = (pe_30_done & (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_30_read_in = (!(par_done_reg81_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg129_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg195_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg273_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg357_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg441_out | left_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? l3_read_data : '0;
  assign left_30_read_write_en = (!(par_done_reg81_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg129_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg195_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg273_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg357_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg441_out | left_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_30_read_in = (!(par_done_reg71_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg114_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg174_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg330_out | top_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg414_out | top_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_20_write_out : '0;
  assign top_30_read_write_en = (!(par_done_reg71_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg114_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg174_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg330_out | top_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg414_out | top_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_30_top = (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_30_read_out : '0;
  assign pe_30_left = (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_30_read_out : '0;
  assign pe_30_go = (!pe_30_done & (!(par_done_reg101_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg156_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg390_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg472_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_25_write_in = (pe_25_done & (!(par_done_reg389_out | down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg471_out | down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg547_out | down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg611_out | down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg659_out | down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg692_out | down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_25_down : '0;
  assign down_25_write_write_en = (pe_25_done & (!(par_done_reg389_out | down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg471_out | down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg547_out | down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg611_out | down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg659_out | down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg692_out | down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_25_read_in = (!(par_done_reg356_out | left_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg440_out | left_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg520_out | left_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg590_out | left_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg644_out | left_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg682_out | left_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_24_write_out : '0;
  assign left_25_read_write_en = (!(par_done_reg356_out | left_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg440_out | left_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg520_out | left_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg590_out | left_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg644_out | left_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg682_out | left_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_25_read_in = (!(par_done_reg329_out | top_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg413_out | top_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg495_out | top_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg569_out | top_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg629_out | top_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg672_out | top_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_15_write_out : '0;
  assign top_25_read_write_en = (!(par_done_reg329_out | top_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg413_out | top_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg495_out | top_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg569_out | top_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg629_out | top_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg672_out | top_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_25_top = (!(par_done_reg389_out | down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg471_out | down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg547_out | down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg611_out | down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg659_out | down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg692_out | down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_25_read_out : '0;
  assign pe_25_left = (!(par_done_reg389_out | down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg471_out | down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg547_out | down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg611_out | down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg659_out | down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg692_out | down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_25_read_out : '0;
  assign pe_25_go = (!pe_25_done & (!(par_done_reg389_out | down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg471_out | down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg547_out | down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg611_out | down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg659_out | down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg692_out | down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_24_write_in = (pe_24_done & (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_24_down : '0;
  assign down_24_write_write_en = (pe_24_done & (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_24_write_in = (pe_24_done & (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_24_right : '0;
  assign right_24_write_write_en = (pe_24_done & (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_24_read_in = (!(par_done_reg272_out | left_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg355_out | left_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg439_out | left_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg519_out | left_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg589_out | left_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg643_out | left_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_23_write_out : '0;
  assign left_24_read_write_en = (!(par_done_reg272_out | left_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg355_out | left_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg439_out | left_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg519_out | left_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg589_out | left_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg643_out | left_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_24_read_in = (!(par_done_reg247_out | top_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg328_out | top_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg412_out | top_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg494_out | top_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg568_out | top_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg628_out | top_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_14_write_out : '0;
  assign top_24_read_write_en = (!(par_done_reg247_out | top_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg328_out | top_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg412_out | top_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg494_out | top_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg568_out | top_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg628_out | top_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_24_top = (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_24_read_out : '0;
  assign pe_24_left = (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_24_read_out : '0;
  assign pe_24_go = (!pe_24_done & (!(par_done_reg305_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg388_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg470_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg546_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg610_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg658_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_23_write_in = (pe_23_done & (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_23_down : '0;
  assign down_23_write_write_en = (pe_23_done & (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_23_write_in = (pe_23_done & (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_23_right : '0;
  assign right_23_write_write_en = (pe_23_done & (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_23_read_in = (!(par_done_reg194_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg271_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg354_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg438_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg518_out | left_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg588_out | left_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_22_write_out : '0;
  assign left_23_read_write_en = (!(par_done_reg194_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg271_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg354_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg438_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg518_out | left_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg588_out | left_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_23_read_in = (!(par_done_reg173_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg246_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg327_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg411_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg493_out | top_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg567_out | top_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_13_write_out : '0;
  assign top_23_read_write_en = (!(par_done_reg173_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg246_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg327_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg411_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg493_out | top_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg567_out | top_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_23_top = (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_23_read_out : '0;
  assign pe_23_left = (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_23_read_out : '0;
  assign pe_23_go = (!pe_23_done & (!(par_done_reg225_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg304_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg387_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg469_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg545_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg609_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_22_write_in = (pe_22_done & (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_22_down : '0;
  assign down_22_write_write_en = (pe_22_done & (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_22_write_in = (pe_22_done & (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_22_right : '0;
  assign right_22_write_write_en = (pe_22_done & (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_22_read_in = (!(par_done_reg128_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg193_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg270_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg353_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg437_out | left_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg517_out | left_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_21_write_out : '0;
  assign left_22_read_write_en = (!(par_done_reg128_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg193_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg270_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg353_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg437_out | left_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg517_out | left_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_22_read_in = (!(par_done_reg113_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg172_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg326_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg410_out | top_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg492_out | top_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_12_write_out : '0;
  assign top_22_read_write_en = (!(par_done_reg113_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg172_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg326_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg410_out | top_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg492_out | top_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_22_top = (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_22_read_out : '0;
  assign pe_22_left = (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_22_read_out : '0;
  assign pe_22_go = (!pe_22_done & (!(par_done_reg155_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg224_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg386_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg468_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg544_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_21_write_in = (pe_21_done & (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_21_down : '0;
  assign down_21_write_write_en = (pe_21_done & (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_21_write_in = (pe_21_done & (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_21_right : '0;
  assign right_21_write_write_en = (pe_21_done & (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_21_read_in = (!(par_done_reg80_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg192_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg269_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg352_out | left_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg436_out | left_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_20_write_out : '0;
  assign left_21_read_write_en = (!(par_done_reg80_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg192_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg269_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg352_out | left_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg436_out | left_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_21_read_in = (!(par_done_reg70_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg112_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg171_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg325_out | top_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg409_out | top_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_11_write_out : '0;
  assign top_21_read_write_en = (!(par_done_reg70_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg112_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg171_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg325_out | top_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg409_out | top_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_21_top = (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_21_read_out : '0;
  assign pe_21_left = (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_21_read_out : '0;
  assign pe_21_go = (!pe_21_done & (!(par_done_reg100_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg385_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg467_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_20_write_in = (pe_20_done & (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_20_down : '0;
  assign down_20_write_write_en = (pe_20_done & (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_20_write_in = (pe_20_done & (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_20_right : '0;
  assign right_20_write_write_en = (pe_20_done & (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_20_read_in = (!(par_done_reg47_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg79_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg126_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg191_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg268_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg351_out | left_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? l2_read_data : '0;
  assign left_20_read_write_en = (!(par_done_reg47_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg79_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg126_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg191_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg268_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg351_out | left_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_20_read_in = (!(par_done_reg41_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg69_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg111_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg170_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg243_out | top_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg324_out | top_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_10_write_out : '0;
  assign top_20_read_write_en = (!(par_done_reg41_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg69_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg111_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg170_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg243_out | top_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg324_out | top_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_20_top = (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_20_read_out : '0;
  assign pe_20_left = (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_20_read_out : '0;
  assign pe_20_go = (!pe_20_done & (!(par_done_reg61_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg99_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg384_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_15_write_in = (pe_15_done & (!(par_done_reg300_out | down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg383_out | down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg466_out | down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg543_out | down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg608_out | down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg657_out | down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_15_down : '0;
  assign down_15_write_write_en = (pe_15_done & (!(par_done_reg300_out | down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg383_out | down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg466_out | down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg543_out | down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg608_out | down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg657_out | down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_15_read_in = (!(par_done_reg267_out | left_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg350_out | left_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg435_out | left_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg516_out | left_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg587_out | left_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg642_out | left_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_14_write_out : '0;
  assign left_15_read_write_en = (!(par_done_reg267_out | left_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg350_out | left_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg435_out | left_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg516_out | left_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg587_out | left_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg642_out | left_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_15_read_in = (!(par_done_reg242_out | top_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg323_out | top_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg408_out | top_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg491_out | top_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg566_out | top_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg627_out | top_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_05_write_out : '0;
  assign top_15_read_write_en = (!(par_done_reg242_out | top_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg323_out | top_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg408_out | top_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg491_out | top_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg566_out | top_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg627_out | top_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_15_top = (!(par_done_reg300_out | down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg383_out | down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg466_out | down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg543_out | down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg608_out | down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg657_out | down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_15_read_out : '0;
  assign pe_15_left = (!(par_done_reg300_out | down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg383_out | down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg466_out | down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg543_out | down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg608_out | down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg657_out | down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_15_read_out : '0;
  assign pe_15_go = (!pe_15_done & (!(par_done_reg300_out | down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg383_out | down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg466_out | down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg543_out | down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg608_out | down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg657_out | down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_14_write_in = (pe_14_done & (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_14_down : '0;
  assign down_14_write_write_en = (pe_14_done & (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_14_write_in = (pe_14_done & (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_14_right : '0;
  assign right_14_write_write_en = (pe_14_done & (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_14_read_in = (!(par_done_reg190_out | left_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg266_out | left_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg349_out | left_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg434_out | left_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg515_out | left_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg586_out | left_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_13_write_out : '0;
  assign left_14_read_write_en = (!(par_done_reg190_out | left_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg266_out | left_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg349_out | left_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg434_out | left_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg515_out | left_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg586_out | left_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_14_read_in = (!(par_done_reg169_out | top_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | top_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg322_out | top_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg407_out | top_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg490_out | top_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg565_out | top_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_04_write_out : '0;
  assign top_14_read_write_en = (!(par_done_reg169_out | top_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | top_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg322_out | top_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg407_out | top_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg490_out | top_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg565_out | top_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_14_top = (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_14_read_out : '0;
  assign pe_14_left = (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_14_read_out : '0;
  assign pe_14_go = (!pe_14_done & (!(par_done_reg221_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg382_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg465_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg542_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg607_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_13_write_in = (pe_13_done & (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_13_down : '0;
  assign down_13_write_write_en = (pe_13_done & (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_13_write_in = (pe_13_done & (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_13_right : '0;
  assign right_13_write_write_en = (pe_13_done & (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_13_read_in = (!(par_done_reg125_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg189_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg265_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg348_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg433_out | left_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg514_out | left_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_12_write_out : '0;
  assign left_13_read_write_en = (!(par_done_reg125_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg189_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg265_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg348_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg433_out | left_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg514_out | left_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_13_read_in = (!(par_done_reg110_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg168_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg321_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg406_out | top_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg489_out | top_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_03_write_out : '0;
  assign top_13_read_write_en = (!(par_done_reg110_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg168_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg321_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg406_out | top_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg489_out | top_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_13_top = (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_13_read_out : '0;
  assign pe_13_left = (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_13_read_out : '0;
  assign pe_13_go = (!pe_13_done & (!(par_done_reg152_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg381_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg464_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg541_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_12_write_in = (pe_12_done & (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_12_down : '0;
  assign down_12_write_write_en = (pe_12_done & (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_12_write_in = (pe_12_done & (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_12_right : '0;
  assign right_12_write_write_en = (pe_12_done & (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_12_read_in = (!(par_done_reg78_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg188_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg264_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg347_out | left_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg432_out | left_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_11_write_out : '0;
  assign left_12_read_write_en = (!(par_done_reg78_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg188_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg264_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg347_out | left_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg432_out | left_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_12_read_in = (!(par_done_reg68_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg239_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg320_out | top_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg405_out | top_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_02_write_out : '0;
  assign top_12_read_write_en = (!(par_done_reg68_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg239_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg320_out | top_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg405_out | top_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_12_top = (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_12_read_out : '0;
  assign pe_12_left = (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_12_read_out : '0;
  assign pe_12_go = (!pe_12_done & (!(par_done_reg98_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg380_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg463_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_11_write_in = (pe_11_done & (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_11_down : '0;
  assign down_11_write_write_en = (pe_11_done & (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_11_write_in = (pe_11_done & (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_11_right : '0;
  assign right_11_write_write_en = (pe_11_done & (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_11_read_in = (!(par_done_reg46_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg123_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg263_out | left_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg346_out | left_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_10_write_out : '0;
  assign left_11_read_write_en = (!(par_done_reg46_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg123_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg263_out | left_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg346_out | left_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_11_read_in = (!(par_done_reg40_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg238_out | top_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg319_out | top_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? down_01_write_out : '0;
  assign top_11_read_write_en = (!(par_done_reg40_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg238_out | top_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg319_out | top_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_11_top = (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_11_read_out : '0;
  assign pe_11_left = (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_11_read_out : '0;
  assign pe_11_go = (!pe_11_done & (!(par_done_reg60_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg218_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg379_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_10_write_in = (pe_10_done & (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_10_down : '0;
  assign down_10_write_write_en = (pe_10_done & (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_10_write_in = (pe_10_done & (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_10_right : '0;
  assign right_10_write_write_en = (pe_10_done & (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_10_read_in = (!(par_done_reg26_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg45_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg76_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg186_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg262_out | left_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? l1_read_data : '0;
  assign left_10_read_write_en = (!(par_done_reg26_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg45_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg76_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg186_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg262_out | left_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_10_read_in = (!(par_done_reg23_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg66_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg165_out | top_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg237_out | top_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? down_00_write_out : '0;
  assign top_10_read_write_en = (!(par_done_reg23_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg39_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg66_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg165_out | top_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg237_out | top_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_10_top = (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_10_read_out : '0;
  assign pe_10_left = (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_10_read_out : '0;
  assign pe_10_go = (!pe_10_done & (!(par_done_reg35_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg59_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg295_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_05_write_in = (pe_05_done & (!(par_done_reg216_out | down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg294_out | down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg378_out | down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg462_out | down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg540_out | down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg606_out | down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_05_down : '0;
  assign down_05_write_write_en = (pe_05_done & (!(par_done_reg216_out | down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg294_out | down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg378_out | down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg462_out | down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg540_out | down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg606_out | down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_05_read_in = (!(par_done_reg185_out | left_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg261_out | left_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg345_out | left_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg431_out | left_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg513_out | left_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg585_out | left_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_04_write_out : '0;
  assign left_05_read_write_en = (!(par_done_reg185_out | left_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg261_out | left_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg345_out | left_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg431_out | left_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg513_out | left_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg585_out | left_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_05_read_in = (!(par_done_reg164_out | top_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg236_out | top_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg318_out | top_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg404_out | top_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg488_out | top_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg564_out | top_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? t5_read_data : '0;
  assign top_05_read_write_en = (!(par_done_reg164_out | top_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg236_out | top_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg318_out | top_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg404_out | top_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg488_out | top_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg564_out | top_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_05_top = (!(par_done_reg216_out | down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg294_out | down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg378_out | down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg462_out | down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg540_out | down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg606_out | down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_05_read_out : '0;
  assign pe_05_left = (!(par_done_reg216_out | down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg294_out | down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg378_out | down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg462_out | down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg540_out | down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg606_out | down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_05_read_out : '0;
  assign pe_05_go = (!pe_05_done & (!(par_done_reg216_out | down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg294_out | down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg378_out | down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg462_out | down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg540_out | down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg606_out | down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_04_write_in = (pe_04_done & (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_04_down : '0;
  assign down_04_write_write_en = (pe_04_done & (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_04_write_in = (pe_04_done & (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_04_right : '0;
  assign right_04_write_write_en = (pe_04_done & (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_04_read_in = (!(par_done_reg121_out | left_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg260_out | left_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg344_out | left_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg430_out | left_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg512_out | left_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_03_write_out : '0;
  assign left_04_read_write_en = (!(par_done_reg121_out | left_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg260_out | left_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg344_out | left_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg430_out | left_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg512_out | left_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_04_read_in = (!(par_done_reg106_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg235_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg317_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg403_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg487_out | top_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? t4_read_data : '0;
  assign top_04_read_write_en = (!(par_done_reg106_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg235_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg317_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg403_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg487_out | top_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_04_top = (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_04_read_out : '0;
  assign pe_04_left = (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_04_read_out : '0;
  assign pe_04_go = (!pe_04_done & (!(par_done_reg148_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg293_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg377_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg461_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg539_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_03_write_in = (pe_03_done & (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_03_down : '0;
  assign down_03_write_write_en = (pe_03_done & (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_03_write_in = (pe_03_done & (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_03_right : '0;
  assign right_03_write_write_en = (pe_03_done & (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_03_read_in = (!(par_done_reg75_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg120_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg183_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg259_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg343_out | left_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg429_out | left_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_02_write_out : '0;
  assign left_03_read_write_en = (!(par_done_reg75_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg120_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg183_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg259_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg343_out | left_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg429_out | left_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_03_read_in = (!(par_done_reg65_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg105_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg162_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg234_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg316_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg402_out | top_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? t3_read_data : '0;
  assign top_03_read_write_en = (!(par_done_reg65_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg105_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg162_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg234_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg316_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg402_out | top_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_03_top = (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_03_read_out : '0;
  assign pe_03_left = (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_03_read_out : '0;
  assign pe_03_go = (!pe_03_done & (!(par_done_reg95_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg147_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg292_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg376_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg460_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_02_write_in = (pe_02_done & (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_02_down : '0;
  assign down_02_write_write_en = (pe_02_done & (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_02_write_in = (pe_02_done & (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_02_right : '0;
  assign right_02_write_write_en = (pe_02_done & (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_02_read_in = (!(par_done_reg44_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg74_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg119_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg182_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg258_out | left_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg342_out | left_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? right_01_write_out : '0;
  assign left_02_read_write_en = (!(par_done_reg44_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg74_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg119_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg182_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg258_out | left_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg342_out | left_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_02_read_in = (!(par_done_reg38_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg104_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg161_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg233_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg315_out | top_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? t2_read_data : '0;
  assign top_02_read_write_en = (!(par_done_reg38_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg104_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg161_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg233_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg315_out | top_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_02_top = (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_02_read_out : '0;
  assign pe_02_left = (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_02_read_out : '0;
  assign pe_02_go = (!pe_02_done & (!(par_done_reg58_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg291_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg375_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign down_01_write_in = (pe_01_done & (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_01_down : '0;
  assign down_01_write_write_en = (pe_01_done & (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign right_01_write_in = (pe_01_done & (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? pe_01_right : '0;
  assign right_01_write_write_en = (pe_01_done & (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign left_01_read_in = (!(par_done_reg25_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg73_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg118_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg181_out | left_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg257_out | left_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? right_00_write_out : '0;
  assign left_01_read_write_en = (!(par_done_reg25_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg73_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg118_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg181_out | left_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg257_out | left_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign top_01_read_in = (!(par_done_reg22_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg63_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg103_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg160_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg232_out | top_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? t1_read_data : '0;
  assign top_01_read_write_en = (!(par_done_reg22_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg63_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg103_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg160_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg232_out | top_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign pe_01_top = (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? top_01_read_out : '0;
  assign pe_01_left = (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? left_01_read_out : '0;
  assign pe_01_go = (!pe_01_done & (!(par_done_reg34_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg212_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg290_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go)) ? 1'd1 : '0;
  assign down_00_write_in = (pe_00_done & (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_00_down : '0;
  assign down_00_write_write_en = (pe_00_done & (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign right_00_write_in = (pe_00_done & (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? pe_00_right : '0;
  assign right_00_write_write_en = (pe_00_done & (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign left_00_read_in = (!(par_done_reg15_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg24_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg42_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg117_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg180_out | left_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? l0_read_data : '0;
  assign left_00_read_write_en = (!(par_done_reg15_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg24_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg42_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg117_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg180_out | left_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign top_00_read_in = (!(par_done_reg14_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg21_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg36_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg159_out | top_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? t0_read_data : '0;
  assign top_00_read_write_en = (!(par_done_reg14_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg21_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg36_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg159_out | top_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign pe_00_top = (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? top_00_read_out : '0;
  assign pe_00_left = (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? left_00_read_out : '0;
  assign pe_00_go = (!pe_00_done & (!(par_done_reg20_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg56_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go)) ? 1'd1 : '0;
  assign l5_addr0 = (!(par_done_reg200_out | left_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg280_out | left_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg366_out | left_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg452_out | left_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg532_out | left_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg600_out | left_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? l5_idx_out : '0;
  assign l5_add_left = (!(par_done_reg143_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg289_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg374_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg459_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg538_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 3'd1 : '0;
  assign l5_add_right = (!(par_done_reg143_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg289_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg374_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg459_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg538_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? l5_idx_out : '0;
  assign l5_idx_in = (!(par_done_reg143_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg289_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg374_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg459_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg538_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? l5_add_out : (!(par_done_reg11_out | l5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l5_idx_write_en = (!(par_done_reg11_out | l5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg143_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg289_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg374_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg459_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg538_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign l4_addr0 = (!(par_done_reg131_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg198_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg277_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg362_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg447_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg526_out | left_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? l4_idx_out : '0;
  assign l4_add_left = (!(par_done_reg91_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg142_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg288_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg373_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg458_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 3'd1 : '0;
  assign l4_add_right = (!(par_done_reg91_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg142_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg288_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg373_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg458_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? l4_idx_out : '0;
  assign l4_idx_in = (!(par_done_reg91_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg142_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg288_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg373_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg458_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? l4_add_out : (!(par_done_reg10_out | l4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l4_idx_write_en = (!(par_done_reg10_out | l4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg91_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg142_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg288_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg373_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg458_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign l3_addr0 = (!(par_done_reg81_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg129_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg195_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg273_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg357_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg441_out | left_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? l3_idx_out : '0;
  assign l3_add_left = (!(par_done_reg55_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg287_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg372_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 3'd1 : '0;
  assign l3_add_right = (!(par_done_reg55_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg287_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg372_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? l3_idx_out : '0;
  assign l3_idx_in = (!(par_done_reg55_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg287_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg372_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? l3_add_out : (!(par_done_reg9_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l3_idx_write_en = (!(par_done_reg9_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg55_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg287_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg372_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign l2_addr0 = (!(par_done_reg47_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg79_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg126_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg191_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg268_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg351_out | left_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? l2_idx_out : '0;
  assign l2_add_left = (!(par_done_reg32_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg286_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 3'd1 : '0;
  assign l2_add_right = (!(par_done_reg32_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg286_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? l2_idx_out : '0;
  assign l2_idx_in = (!(par_done_reg32_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg286_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? l2_add_out : (!(par_done_reg8_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l2_idx_write_en = (!(par_done_reg8_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg32_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg286_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign l1_addr0 = (!(par_done_reg26_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg45_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg76_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg186_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg262_out | left_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? l1_idx_out : '0;
  assign l1_add_left = (!(par_done_reg19_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 3'd1 : '0;
  assign l1_add_right = (!(par_done_reg19_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? l1_idx_out : '0;
  assign l1_idx_in = (!(par_done_reg19_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? l1_add_out : (!(par_done_reg7_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l1_idx_write_en = (!(par_done_reg7_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg19_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign l0_addr0 = (!(par_done_reg15_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg24_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg42_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg72_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg117_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg180_out | left_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? l0_idx_out : '0;
  assign l0_add_left = (!(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg28_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 3'd1 : '0;
  assign l0_add_right = (!(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg28_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? l0_idx_out : '0;
  assign l0_idx_in = (!(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg28_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? l0_add_out : (!(par_done_reg6_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign l0_idx_write_en = (!(par_done_reg6_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg13_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg28_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg49_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg83_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg133_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign t5_addr0 = (!(par_done_reg164_out | top_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg236_out | top_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg318_out | top_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg404_out | top_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg488_out | top_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg564_out | top_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? t5_idx_out : '0;
  assign t5_add_left = (!(par_done_reg138_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg285_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg371_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg457_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg537_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 3'd1 : '0;
  assign t5_add_right = (!(par_done_reg138_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg285_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg371_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg457_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg537_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? t5_idx_out : '0;
  assign t5_idx_in = (!(par_done_reg138_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg285_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg371_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg457_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg537_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? t5_add_out : (!(par_done_reg5_out | t5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t5_idx_write_en = (!(par_done_reg5_out | t5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg138_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg285_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg371_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg457_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg537_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign t4_addr0 = (!(par_done_reg106_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg235_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg317_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg403_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg487_out | top_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? t4_idx_out : '0;
  assign t4_add_left = (!(par_done_reg87_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg284_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg370_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg456_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 3'd1 : '0;
  assign t4_add_right = (!(par_done_reg87_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg284_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg370_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg456_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? t4_idx_out : '0;
  assign t4_idx_in = (!(par_done_reg87_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg284_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg370_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg456_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? t4_add_out : (!(par_done_reg4_out | t4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t4_idx_write_en = (!(par_done_reg4_out | t4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg87_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg204_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg284_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg370_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg456_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign t3_addr0 = (!(par_done_reg65_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg105_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg162_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg234_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg316_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg402_out | top_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? t3_idx_out : '0;
  assign t3_add_left = (!(par_done_reg52_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg203_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg283_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg369_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 3'd1 : '0;
  assign t3_add_right = (!(par_done_reg52_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg203_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg283_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg369_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? t3_idx_out : '0;
  assign t3_idx_in = (!(par_done_reg52_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg203_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg283_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg369_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? t3_add_out : (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t3_idx_write_en = (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg52_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg203_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg283_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg369_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign t2_addr0 = (!(par_done_reg38_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg64_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg104_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg161_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg233_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg315_out | top_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? t2_idx_out : '0;
  assign t2_add_left = (!(par_done_reg30_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg282_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 3'd1 : '0;
  assign t2_add_right = (!(par_done_reg30_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg282_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? t2_idx_out : '0;
  assign t2_idx_in = (!(par_done_reg30_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg282_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? t2_add_out : (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t2_idx_write_en = (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg30_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg51_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg85_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg135_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg202_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg282_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign t1_addr0 = (!(par_done_reg22_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg37_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg63_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg103_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg160_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg232_out | top_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go) ? t1_idx_out : '0;
  assign t1_add_left = (!(par_done_reg18_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 3'd1 : '0;
  assign t1_add_right = (!(par_done_reg18_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? t1_idx_out : '0;
  assign t1_idx_in = (!(par_done_reg18_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? t1_add_out : (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t1_idx_write_en = (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg18_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg29_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg50_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg84_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg134_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg201_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign t0_addr0 = (!(par_done_reg14_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg21_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg36_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg62_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg102_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg159_out | top_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go) ? t0_idx_out : '0;
  assign t0_add_left = (!(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 3'd1 : '0;
  assign t0_add_right = (!(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? t0_idx_out : '0;
  assign t0_idx_in = (!(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? t0_add_out : (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 3'd7 : '0;
  assign t0_idx_write_en = (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg12_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg27_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg48_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg82_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg132_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_reset0_in = par_reset0_out ? 1'd0 : (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & par_done_reg8_out & par_done_reg9_out & par_done_reg10_out & par_done_reg11_out & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_reset0_write_en = (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & par_done_reg8_out & par_done_reg9_out & par_done_reg10_out & par_done_reg11_out & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg0_in = par_reset0_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg0_write_en = (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg1_in = par_reset0_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg1_write_en = (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg2_in = par_reset0_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg2_write_en = (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg3_in = par_reset0_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg3_write_en = (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg4_in = par_reset0_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg4_write_en = (t4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg5_in = par_reset0_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg5_write_en = (t5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg6_in = par_reset0_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg6_write_en = (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg7_in = par_reset0_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg7_write_en = (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg8_in = par_reset0_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg8_write_en = (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg9_in = par_reset0_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg9_write_en = (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg10_in = par_reset0_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg10_write_en = (l4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg11_in = par_reset0_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg11_write_en = (l5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_reset1_in = par_reset1_out ? 1'd0 : (par_done_reg12_out & par_done_reg13_out & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_reset1_write_en = (par_done_reg12_out & par_done_reg13_out & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg12_in = par_reset1_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg12_write_en = (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg13_in = par_reset1_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg13_write_en = (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_reset2_in = par_reset2_out ? 1'd0 : (par_done_reg14_out & par_done_reg15_out & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_reset2_write_en = (par_done_reg14_out & par_done_reg15_out & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg14_in = par_reset2_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg14_write_en = (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg15_in = par_reset2_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg15_write_en = (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_reset3_in = par_reset3_out ? 1'd0 : (par_done_reg16_out & par_done_reg17_out & par_done_reg18_out & par_done_reg19_out & par_done_reg20_out & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_reset3_write_en = (par_done_reg16_out & par_done_reg17_out & par_done_reg18_out & par_done_reg19_out & par_done_reg20_out & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg16_in = par_reset3_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg16_write_en = (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg17_in = par_reset3_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg17_write_en = (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg18_in = par_reset3_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg18_write_en = (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg19_in = par_reset3_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg19_write_en = (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg20_in = par_reset3_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg20_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_reset4_in = par_reset4_out ? 1'd0 : (par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & par_done_reg25_out & par_done_reg26_out & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_reset4_write_en = (par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & par_done_reg25_out & par_done_reg26_out & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg21_in = par_reset4_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg21_write_en = (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg22_in = par_reset4_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg22_write_en = (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg23_in = par_reset4_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg23_write_en = (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg24_in = par_reset4_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg24_write_en = (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg25_in = par_reset4_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg25_write_en = (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg26_in = par_reset4_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg26_write_en = (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_reset5_in = par_reset5_out ? 1'd0 : (par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_reset5_write_en = (par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg27_in = par_reset5_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg27_write_en = (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg28_in = par_reset5_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg28_write_en = (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg29_in = par_reset5_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg29_write_en = (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg30_in = par_reset5_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg30_write_en = (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg31_in = par_reset5_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg31_write_en = (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg32_in = par_reset5_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg32_write_en = (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg33_in = par_reset5_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg33_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg34_in = par_reset5_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg34_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg35_in = par_reset5_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg35_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_reset6_in = par_reset6_out ? 1'd0 : (par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_reset6_write_en = (par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg36_in = par_reset6_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg36_write_en = (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg37_in = par_reset6_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg37_write_en = (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg38_in = par_reset6_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg38_write_en = (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg39_in = par_reset6_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg39_write_en = (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg40_in = par_reset6_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg40_write_en = (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg41_in = par_reset6_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg41_write_en = (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg42_in = par_reset6_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg42_write_en = (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg43_in = par_reset6_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg43_write_en = (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg44_in = par_reset6_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg44_write_en = (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg45_in = par_reset6_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg45_write_en = (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg46_in = par_reset6_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg46_write_en = (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg47_in = par_reset6_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg47_write_en = (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_reset7_in = par_reset7_out ? 1'd0 : (par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_reset7_write_en = (par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg48_in = par_reset7_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg48_write_en = (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg49_in = par_reset7_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg49_write_en = (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg50_in = par_reset7_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg50_write_en = (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg51_in = par_reset7_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg51_write_en = (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg52_in = par_reset7_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg52_write_en = (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg53_in = par_reset7_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg53_write_en = (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg54_in = par_reset7_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg54_write_en = (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg55_in = par_reset7_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg55_write_en = (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg56_in = par_reset7_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg56_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg57_in = par_reset7_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg57_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg58_in = par_reset7_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg58_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg59_in = par_reset7_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg59_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg60_in = par_reset7_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg60_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg61_in = par_reset7_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg61_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_reset8_in = par_reset8_out ? 1'd0 : (par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_reset8_write_en = (par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg62_in = par_reset8_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg62_write_en = (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg63_in = par_reset8_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg63_write_en = (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg64_in = par_reset8_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg64_write_en = (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg65_in = par_reset8_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg65_write_en = (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg66_in = par_reset8_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg66_write_en = (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg67_in = par_reset8_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg67_write_en = (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg68_in = par_reset8_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg68_write_en = (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg69_in = par_reset8_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg69_write_en = (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg70_in = par_reset8_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg70_write_en = (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg71_in = par_reset8_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg71_write_en = (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg72_in = par_reset8_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg72_write_en = (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg73_in = par_reset8_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg73_write_en = (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg74_in = par_reset8_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg74_write_en = (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg75_in = par_reset8_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg75_write_en = (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg76_in = par_reset8_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg76_write_en = (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg77_in = par_reset8_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg77_write_en = (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg78_in = par_reset8_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg78_write_en = (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg79_in = par_reset8_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg79_write_en = (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg80_in = par_reset8_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg80_write_en = (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg81_in = par_reset8_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg81_write_en = (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_reset9_in = par_reset9_out ? 1'd0 : (par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_reset9_write_en = (par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg82_in = par_reset9_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg82_write_en = (t0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg83_in = par_reset9_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg83_write_en = (l0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg84_in = par_reset9_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg84_write_en = (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg85_in = par_reset9_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg85_write_en = (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg86_in = par_reset9_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg86_write_en = (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg87_in = par_reset9_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg87_write_en = (t4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg88_in = par_reset9_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg88_write_en = (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg89_in = par_reset9_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg89_write_en = (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg90_in = par_reset9_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg90_write_en = (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg91_in = par_reset9_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg91_write_en = (l4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg92_in = par_reset9_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg92_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg93_in = par_reset9_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg93_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg94_in = par_reset9_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg94_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg95_in = par_reset9_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg95_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg96_in = par_reset9_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg96_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg97_in = par_reset9_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg97_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg98_in = par_reset9_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg98_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg99_in = par_reset9_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg99_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg100_in = par_reset9_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg100_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg101_in = par_reset9_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg101_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_reset10_in = par_reset10_out ? 1'd0 : (par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & par_done_reg130_out & par_done_reg131_out & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_reset10_write_en = (par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & par_done_reg130_out & par_done_reg131_out & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg102_in = par_reset10_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg102_write_en = (top_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg103_in = par_reset10_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg103_write_en = (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg104_in = par_reset10_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg104_write_en = (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg105_in = par_reset10_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg105_write_en = (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg106_in = par_reset10_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg106_write_en = (top_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg107_in = par_reset10_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg107_write_en = (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg108_in = par_reset10_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg108_write_en = (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg109_in = par_reset10_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg109_write_en = (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg110_in = par_reset10_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg110_write_en = (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg111_in = par_reset10_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg111_write_en = (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg112_in = par_reset10_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg112_write_en = (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg113_in = par_reset10_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg113_write_en = (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg114_in = par_reset10_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg114_write_en = (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg115_in = par_reset10_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg115_write_en = (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg116_in = par_reset10_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg116_write_en = (top_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg117_in = par_reset10_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg117_write_en = (left_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg118_in = par_reset10_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg118_write_en = (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg119_in = par_reset10_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg119_write_en = (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg120_in = par_reset10_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg120_write_en = (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg121_in = par_reset10_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg121_write_en = (left_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg122_in = par_reset10_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg122_write_en = (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg123_in = par_reset10_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg123_write_en = (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg124_in = par_reset10_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg124_write_en = (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg125_in = par_reset10_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg125_write_en = (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg126_in = par_reset10_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg126_write_en = (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg127_in = par_reset10_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg127_write_en = (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg128_in = par_reset10_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg128_write_en = (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg129_in = par_reset10_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg129_write_en = (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg130_in = par_reset10_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg130_write_en = (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg131_in = par_reset10_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg131_write_en = (left_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_reset11_in = par_reset11_out ? 1'd0 : (par_done_reg132_out & par_done_reg133_out & par_done_reg134_out & par_done_reg135_out & par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & par_done_reg158_out & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_reset11_write_en = (par_done_reg132_out & par_done_reg133_out & par_done_reg134_out & par_done_reg135_out & par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & par_done_reg158_out & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg132_in = par_reset11_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg132_write_en = (t0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg133_in = par_reset11_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg133_write_en = (l0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg134_in = par_reset11_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg134_write_en = (t1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg135_in = par_reset11_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg135_write_en = (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg136_in = par_reset11_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg136_write_en = (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg137_in = par_reset11_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg137_write_en = (t4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg138_in = par_reset11_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg138_write_en = (t5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg139_in = par_reset11_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg139_write_en = (l1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg140_in = par_reset11_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg140_write_en = (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg141_in = par_reset11_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg141_write_en = (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg142_in = par_reset11_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg142_write_en = (l4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg143_in = par_reset11_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg143_write_en = (l5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg144_in = par_reset11_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg144_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg145_in = par_reset11_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg145_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg146_in = par_reset11_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg146_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg147_in = par_reset11_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg147_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg148_in = par_reset11_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg148_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg149_in = par_reset11_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg149_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg150_in = par_reset11_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg150_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg151_in = par_reset11_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg151_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg152_in = par_reset11_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg152_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg153_in = par_reset11_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg153_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg154_in = par_reset11_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg154_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg155_in = par_reset11_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg155_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg156_in = par_reset11_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg156_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg157_in = par_reset11_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg157_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg158_in = par_reset11_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg158_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_reset12_in = par_reset12_out ? 1'd0 : (par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_reset12_write_en = (par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg159_in = par_reset12_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg159_write_en = (top_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg160_in = par_reset12_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg160_write_en = (top_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg161_in = par_reset12_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg161_write_en = (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg162_in = par_reset12_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg162_write_en = (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg163_in = par_reset12_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg163_write_en = (top_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg164_in = par_reset12_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg164_write_en = (top_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg165_in = par_reset12_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg165_write_en = (top_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg166_in = par_reset12_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg166_write_en = (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg167_in = par_reset12_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg167_write_en = (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg168_in = par_reset12_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg168_write_en = (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg169_in = par_reset12_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg169_write_en = (top_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg170_in = par_reset12_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg170_write_en = (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg171_in = par_reset12_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg171_write_en = (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg172_in = par_reset12_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg172_write_en = (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg173_in = par_reset12_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg173_write_en = (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg174_in = par_reset12_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg174_write_en = (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg175_in = par_reset12_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg175_write_en = (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg176_in = par_reset12_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg176_write_en = (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg177_in = par_reset12_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg177_write_en = (top_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg178_in = par_reset12_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg178_write_en = (top_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg179_in = par_reset12_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg179_write_en = (top_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg180_in = par_reset12_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg180_write_en = (left_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg181_in = par_reset12_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg181_write_en = (left_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg182_in = par_reset12_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg182_write_en = (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg183_in = par_reset12_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg183_write_en = (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg184_in = par_reset12_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg184_write_en = (left_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg185_in = par_reset12_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg185_write_en = (left_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg186_in = par_reset12_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg186_write_en = (left_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg187_in = par_reset12_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg187_write_en = (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg188_in = par_reset12_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg188_write_en = (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg189_in = par_reset12_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg189_write_en = (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg190_in = par_reset12_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg190_write_en = (left_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg191_in = par_reset12_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg191_write_en = (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg192_in = par_reset12_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg192_write_en = (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg193_in = par_reset12_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg193_write_en = (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg194_in = par_reset12_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg194_write_en = (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg195_in = par_reset12_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg195_write_en = (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg196_in = par_reset12_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg196_write_en = (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg197_in = par_reset12_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg197_write_en = (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg198_in = par_reset12_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg198_write_en = (left_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg199_in = par_reset12_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg199_write_en = (left_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg200_in = par_reset12_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg200_write_en = (left_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_reset13_in = par_reset13_out ? 1'd0 : (par_done_reg201_out & par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & par_done_reg213_out & par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & par_done_reg229_out & par_done_reg230_out & par_done_reg231_out & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_reset13_write_en = (par_done_reg201_out & par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & par_done_reg213_out & par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & par_done_reg229_out & par_done_reg230_out & par_done_reg231_out & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg201_in = par_reset13_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg201_write_en = (t1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg202_in = par_reset13_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg202_write_en = (t2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg203_in = par_reset13_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg203_write_en = (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg204_in = par_reset13_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg204_write_en = (t4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg205_in = par_reset13_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg205_write_en = (t5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg206_in = par_reset13_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg206_write_en = (l1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg207_in = par_reset13_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg207_write_en = (l2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg208_in = par_reset13_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg208_write_en = (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg209_in = par_reset13_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg209_write_en = (l4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg210_in = par_reset13_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg210_write_en = (l5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg211_in = par_reset13_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg211_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg212_in = par_reset13_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg212_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg213_in = par_reset13_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg213_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg214_in = par_reset13_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg214_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg215_in = par_reset13_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg215_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg216_in = par_reset13_out ? 1'd0 : (down_05_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg216_write_en = (down_05_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg217_in = par_reset13_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg217_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg218_in = par_reset13_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg218_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg219_in = par_reset13_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg219_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg220_in = par_reset13_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg220_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg221_in = par_reset13_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg221_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg222_in = par_reset13_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg222_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg223_in = par_reset13_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg223_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg224_in = par_reset13_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg224_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg225_in = par_reset13_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg225_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg226_in = par_reset13_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg226_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg227_in = par_reset13_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg227_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg228_in = par_reset13_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg228_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg229_in = par_reset13_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg229_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg230_in = par_reset13_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg230_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg231_in = par_reset13_out ? 1'd0 : (right_50_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg231_write_en = (right_50_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_reset14_in = par_reset14_out ? 1'd0 : (par_done_reg232_out & par_done_reg233_out & par_done_reg234_out & par_done_reg235_out & par_done_reg236_out & par_done_reg237_out & par_done_reg238_out & par_done_reg239_out & par_done_reg240_out & par_done_reg241_out & par_done_reg242_out & par_done_reg243_out & par_done_reg244_out & par_done_reg245_out & par_done_reg246_out & par_done_reg247_out & par_done_reg248_out & par_done_reg249_out & par_done_reg250_out & par_done_reg251_out & par_done_reg252_out & par_done_reg253_out & par_done_reg254_out & par_done_reg255_out & par_done_reg256_out & par_done_reg257_out & par_done_reg258_out & par_done_reg259_out & par_done_reg260_out & par_done_reg261_out & par_done_reg262_out & par_done_reg263_out & par_done_reg264_out & par_done_reg265_out & par_done_reg266_out & par_done_reg267_out & par_done_reg268_out & par_done_reg269_out & par_done_reg270_out & par_done_reg271_out & par_done_reg272_out & par_done_reg273_out & par_done_reg274_out & par_done_reg275_out & par_done_reg276_out & par_done_reg277_out & par_done_reg278_out & par_done_reg279_out & par_done_reg280_out & par_done_reg281_out & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_reset14_write_en = (par_done_reg232_out & par_done_reg233_out & par_done_reg234_out & par_done_reg235_out & par_done_reg236_out & par_done_reg237_out & par_done_reg238_out & par_done_reg239_out & par_done_reg240_out & par_done_reg241_out & par_done_reg242_out & par_done_reg243_out & par_done_reg244_out & par_done_reg245_out & par_done_reg246_out & par_done_reg247_out & par_done_reg248_out & par_done_reg249_out & par_done_reg250_out & par_done_reg251_out & par_done_reg252_out & par_done_reg253_out & par_done_reg254_out & par_done_reg255_out & par_done_reg256_out & par_done_reg257_out & par_done_reg258_out & par_done_reg259_out & par_done_reg260_out & par_done_reg261_out & par_done_reg262_out & par_done_reg263_out & par_done_reg264_out & par_done_reg265_out & par_done_reg266_out & par_done_reg267_out & par_done_reg268_out & par_done_reg269_out & par_done_reg270_out & par_done_reg271_out & par_done_reg272_out & par_done_reg273_out & par_done_reg274_out & par_done_reg275_out & par_done_reg276_out & par_done_reg277_out & par_done_reg278_out & par_done_reg279_out & par_done_reg280_out & par_done_reg281_out & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg232_in = par_reset14_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg232_write_en = (top_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg233_in = par_reset14_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg233_write_en = (top_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg234_in = par_reset14_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg234_write_en = (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg235_in = par_reset14_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg235_write_en = (top_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg236_in = par_reset14_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg236_write_en = (top_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg237_in = par_reset14_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg237_write_en = (top_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg238_in = par_reset14_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg238_write_en = (top_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg239_in = par_reset14_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg239_write_en = (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg240_in = par_reset14_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg240_write_en = (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg241_in = par_reset14_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg241_write_en = (top_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg242_in = par_reset14_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg242_write_en = (top_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg243_in = par_reset14_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg243_write_en = (top_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg244_in = par_reset14_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg244_write_en = (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg245_in = par_reset14_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg245_write_en = (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg246_in = par_reset14_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg246_write_en = (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg247_in = par_reset14_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg247_write_en = (top_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg248_in = par_reset14_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg248_write_en = (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg249_in = par_reset14_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg249_write_en = (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg250_in = par_reset14_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg250_write_en = (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg251_in = par_reset14_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg251_write_en = (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg252_in = par_reset14_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg252_write_en = (top_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg253_in = par_reset14_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg253_write_en = (top_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg254_in = par_reset14_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg254_write_en = (top_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg255_in = par_reset14_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg255_write_en = (top_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg256_in = par_reset14_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg256_write_en = (top_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg257_in = par_reset14_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg257_write_en = (left_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg258_in = par_reset14_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg258_write_en = (left_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg259_in = par_reset14_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg259_write_en = (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg260_in = par_reset14_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg260_write_en = (left_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg261_in = par_reset14_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg261_write_en = (left_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg262_in = par_reset14_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg262_write_en = (left_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg263_in = par_reset14_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg263_write_en = (left_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg264_in = par_reset14_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg264_write_en = (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg265_in = par_reset14_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg265_write_en = (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg266_in = par_reset14_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg266_write_en = (left_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg267_in = par_reset14_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg267_write_en = (left_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg268_in = par_reset14_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg268_write_en = (left_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg269_in = par_reset14_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg269_write_en = (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg270_in = par_reset14_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg270_write_en = (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg271_in = par_reset14_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg271_write_en = (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg272_in = par_reset14_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg272_write_en = (left_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg273_in = par_reset14_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg273_write_en = (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg274_in = par_reset14_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg274_write_en = (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg275_in = par_reset14_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg275_write_en = (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg276_in = par_reset14_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg276_write_en = (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg277_in = par_reset14_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg277_write_en = (left_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg278_in = par_reset14_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg278_write_en = (left_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg279_in = par_reset14_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg279_write_en = (left_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg280_in = par_reset14_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg280_write_en = (left_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg281_in = par_reset14_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg281_write_en = (left_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_reset15_in = par_reset15_out ? 1'd0 : (par_done_reg282_out & par_done_reg283_out & par_done_reg284_out & par_done_reg285_out & par_done_reg286_out & par_done_reg287_out & par_done_reg288_out & par_done_reg289_out & par_done_reg290_out & par_done_reg291_out & par_done_reg292_out & par_done_reg293_out & par_done_reg294_out & par_done_reg295_out & par_done_reg296_out & par_done_reg297_out & par_done_reg298_out & par_done_reg299_out & par_done_reg300_out & par_done_reg301_out & par_done_reg302_out & par_done_reg303_out & par_done_reg304_out & par_done_reg305_out & par_done_reg306_out & par_done_reg307_out & par_done_reg308_out & par_done_reg309_out & par_done_reg310_out & par_done_reg311_out & par_done_reg312_out & par_done_reg313_out & par_done_reg314_out & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_reset15_write_en = (par_done_reg282_out & par_done_reg283_out & par_done_reg284_out & par_done_reg285_out & par_done_reg286_out & par_done_reg287_out & par_done_reg288_out & par_done_reg289_out & par_done_reg290_out & par_done_reg291_out & par_done_reg292_out & par_done_reg293_out & par_done_reg294_out & par_done_reg295_out & par_done_reg296_out & par_done_reg297_out & par_done_reg298_out & par_done_reg299_out & par_done_reg300_out & par_done_reg301_out & par_done_reg302_out & par_done_reg303_out & par_done_reg304_out & par_done_reg305_out & par_done_reg306_out & par_done_reg307_out & par_done_reg308_out & par_done_reg309_out & par_done_reg310_out & par_done_reg311_out & par_done_reg312_out & par_done_reg313_out & par_done_reg314_out & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg282_in = par_reset15_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg282_write_en = (t2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg283_in = par_reset15_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg283_write_en = (t3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg284_in = par_reset15_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg284_write_en = (t4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg285_in = par_reset15_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg285_write_en = (t5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg286_in = par_reset15_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg286_write_en = (l2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg287_in = par_reset15_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg287_write_en = (l3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg288_in = par_reset15_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg288_write_en = (l4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg289_in = par_reset15_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg289_write_en = (l5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg290_in = par_reset15_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg290_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg291_in = par_reset15_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg291_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg292_in = par_reset15_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg292_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg293_in = par_reset15_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg293_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg294_in = par_reset15_out ? 1'd0 : (down_05_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg294_write_en = (down_05_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg295_in = par_reset15_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg295_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg296_in = par_reset15_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg296_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg297_in = par_reset15_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg297_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg298_in = par_reset15_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg298_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg299_in = par_reset15_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg299_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg300_in = par_reset15_out ? 1'd0 : (down_15_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg300_write_en = (down_15_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg301_in = par_reset15_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg301_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg302_in = par_reset15_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg302_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg303_in = par_reset15_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg303_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg304_in = par_reset15_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg304_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg305_in = par_reset15_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg305_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg306_in = par_reset15_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg306_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg307_in = par_reset15_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg307_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg308_in = par_reset15_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg308_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg309_in = par_reset15_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg309_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg310_in = par_reset15_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg310_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg311_in = par_reset15_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg311_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg312_in = par_reset15_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg312_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg313_in = par_reset15_out ? 1'd0 : (right_50_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg313_write_en = (right_50_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg314_in = par_reset15_out ? 1'd0 : (right_51_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg314_write_en = (right_51_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_reset16_in = par_reset16_out ? 1'd0 : (par_done_reg315_out & par_done_reg316_out & par_done_reg317_out & par_done_reg318_out & par_done_reg319_out & par_done_reg320_out & par_done_reg321_out & par_done_reg322_out & par_done_reg323_out & par_done_reg324_out & par_done_reg325_out & par_done_reg326_out & par_done_reg327_out & par_done_reg328_out & par_done_reg329_out & par_done_reg330_out & par_done_reg331_out & par_done_reg332_out & par_done_reg333_out & par_done_reg334_out & par_done_reg335_out & par_done_reg336_out & par_done_reg337_out & par_done_reg338_out & par_done_reg339_out & par_done_reg340_out & par_done_reg341_out & par_done_reg342_out & par_done_reg343_out & par_done_reg344_out & par_done_reg345_out & par_done_reg346_out & par_done_reg347_out & par_done_reg348_out & par_done_reg349_out & par_done_reg350_out & par_done_reg351_out & par_done_reg352_out & par_done_reg353_out & par_done_reg354_out & par_done_reg355_out & par_done_reg356_out & par_done_reg357_out & par_done_reg358_out & par_done_reg359_out & par_done_reg360_out & par_done_reg361_out & par_done_reg362_out & par_done_reg363_out & par_done_reg364_out & par_done_reg365_out & par_done_reg366_out & par_done_reg367_out & par_done_reg368_out & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_reset16_write_en = (par_done_reg315_out & par_done_reg316_out & par_done_reg317_out & par_done_reg318_out & par_done_reg319_out & par_done_reg320_out & par_done_reg321_out & par_done_reg322_out & par_done_reg323_out & par_done_reg324_out & par_done_reg325_out & par_done_reg326_out & par_done_reg327_out & par_done_reg328_out & par_done_reg329_out & par_done_reg330_out & par_done_reg331_out & par_done_reg332_out & par_done_reg333_out & par_done_reg334_out & par_done_reg335_out & par_done_reg336_out & par_done_reg337_out & par_done_reg338_out & par_done_reg339_out & par_done_reg340_out & par_done_reg341_out & par_done_reg342_out & par_done_reg343_out & par_done_reg344_out & par_done_reg345_out & par_done_reg346_out & par_done_reg347_out & par_done_reg348_out & par_done_reg349_out & par_done_reg350_out & par_done_reg351_out & par_done_reg352_out & par_done_reg353_out & par_done_reg354_out & par_done_reg355_out & par_done_reg356_out & par_done_reg357_out & par_done_reg358_out & par_done_reg359_out & par_done_reg360_out & par_done_reg361_out & par_done_reg362_out & par_done_reg363_out & par_done_reg364_out & par_done_reg365_out & par_done_reg366_out & par_done_reg367_out & par_done_reg368_out & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg315_in = par_reset16_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg315_write_en = (top_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg316_in = par_reset16_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg316_write_en = (top_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg317_in = par_reset16_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg317_write_en = (top_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg318_in = par_reset16_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg318_write_en = (top_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg319_in = par_reset16_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg319_write_en = (top_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg320_in = par_reset16_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg320_write_en = (top_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg321_in = par_reset16_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg321_write_en = (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg322_in = par_reset16_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg322_write_en = (top_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg323_in = par_reset16_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg323_write_en = (top_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg324_in = par_reset16_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg324_write_en = (top_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg325_in = par_reset16_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg325_write_en = (top_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg326_in = par_reset16_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg326_write_en = (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg327_in = par_reset16_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg327_write_en = (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg328_in = par_reset16_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg328_write_en = (top_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg329_in = par_reset16_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg329_write_en = (top_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg330_in = par_reset16_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg330_write_en = (top_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg331_in = par_reset16_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg331_write_en = (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg332_in = par_reset16_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg332_write_en = (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg333_in = par_reset16_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg333_write_en = (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg334_in = par_reset16_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg334_write_en = (top_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg335_in = par_reset16_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg335_write_en = (top_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg336_in = par_reset16_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg336_write_en = (top_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg337_in = par_reset16_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg337_write_en = (top_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg338_in = par_reset16_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg338_write_en = (top_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg339_in = par_reset16_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg339_write_en = (top_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg340_in = par_reset16_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg340_write_en = (top_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg341_in = par_reset16_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg341_write_en = (top_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg342_in = par_reset16_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg342_write_en = (left_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg343_in = par_reset16_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg343_write_en = (left_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg344_in = par_reset16_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg344_write_en = (left_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg345_in = par_reset16_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg345_write_en = (left_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg346_in = par_reset16_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg346_write_en = (left_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg347_in = par_reset16_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg347_write_en = (left_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg348_in = par_reset16_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg348_write_en = (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg349_in = par_reset16_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg349_write_en = (left_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg350_in = par_reset16_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg350_write_en = (left_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg351_in = par_reset16_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg351_write_en = (left_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg352_in = par_reset16_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg352_write_en = (left_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg353_in = par_reset16_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg353_write_en = (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg354_in = par_reset16_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg354_write_en = (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg355_in = par_reset16_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg355_write_en = (left_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg356_in = par_reset16_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg356_write_en = (left_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg357_in = par_reset16_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg357_write_en = (left_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg358_in = par_reset16_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg358_write_en = (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg359_in = par_reset16_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg359_write_en = (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg360_in = par_reset16_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg360_write_en = (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg361_in = par_reset16_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg361_write_en = (left_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg362_in = par_reset16_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg362_write_en = (left_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg363_in = par_reset16_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg363_write_en = (left_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg364_in = par_reset16_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg364_write_en = (left_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg365_in = par_reset16_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg365_write_en = (left_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg366_in = par_reset16_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg366_write_en = (left_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg367_in = par_reset16_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg367_write_en = (left_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg368_in = par_reset16_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg368_write_en = (left_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_reset17_in = par_reset17_out ? 1'd0 : (par_done_reg369_out & par_done_reg370_out & par_done_reg371_out & par_done_reg372_out & par_done_reg373_out & par_done_reg374_out & par_done_reg375_out & par_done_reg376_out & par_done_reg377_out & par_done_reg378_out & par_done_reg379_out & par_done_reg380_out & par_done_reg381_out & par_done_reg382_out & par_done_reg383_out & par_done_reg384_out & par_done_reg385_out & par_done_reg386_out & par_done_reg387_out & par_done_reg388_out & par_done_reg389_out & par_done_reg390_out & par_done_reg391_out & par_done_reg392_out & par_done_reg393_out & par_done_reg394_out & par_done_reg395_out & par_done_reg396_out & par_done_reg397_out & par_done_reg398_out & par_done_reg399_out & par_done_reg400_out & par_done_reg401_out & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_reset17_write_en = (par_done_reg369_out & par_done_reg370_out & par_done_reg371_out & par_done_reg372_out & par_done_reg373_out & par_done_reg374_out & par_done_reg375_out & par_done_reg376_out & par_done_reg377_out & par_done_reg378_out & par_done_reg379_out & par_done_reg380_out & par_done_reg381_out & par_done_reg382_out & par_done_reg383_out & par_done_reg384_out & par_done_reg385_out & par_done_reg386_out & par_done_reg387_out & par_done_reg388_out & par_done_reg389_out & par_done_reg390_out & par_done_reg391_out & par_done_reg392_out & par_done_reg393_out & par_done_reg394_out & par_done_reg395_out & par_done_reg396_out & par_done_reg397_out & par_done_reg398_out & par_done_reg399_out & par_done_reg400_out & par_done_reg401_out & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg369_in = par_reset17_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg369_write_en = (t3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg370_in = par_reset17_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg370_write_en = (t4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg371_in = par_reset17_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg371_write_en = (t5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg372_in = par_reset17_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg372_write_en = (l3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg373_in = par_reset17_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg373_write_en = (l4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg374_in = par_reset17_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg374_write_en = (l5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg375_in = par_reset17_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg375_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg376_in = par_reset17_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg376_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg377_in = par_reset17_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg377_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg378_in = par_reset17_out ? 1'd0 : (down_05_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg378_write_en = (down_05_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg379_in = par_reset17_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg379_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg380_in = par_reset17_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg380_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg381_in = par_reset17_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg381_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg382_in = par_reset17_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg382_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg383_in = par_reset17_out ? 1'd0 : (down_15_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg383_write_en = (down_15_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg384_in = par_reset17_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg384_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg385_in = par_reset17_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg385_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg386_in = par_reset17_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg386_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg387_in = par_reset17_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg387_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg388_in = par_reset17_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg388_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg389_in = par_reset17_out ? 1'd0 : (down_25_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg389_write_en = (down_25_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg390_in = par_reset17_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg390_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg391_in = par_reset17_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg391_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg392_in = par_reset17_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg392_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg393_in = par_reset17_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg393_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg394_in = par_reset17_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg394_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg395_in = par_reset17_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg395_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg396_in = par_reset17_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg396_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg397_in = par_reset17_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg397_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg398_in = par_reset17_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg398_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg399_in = par_reset17_out ? 1'd0 : (right_50_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg399_write_en = (right_50_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg400_in = par_reset17_out ? 1'd0 : (right_51_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg400_write_en = (right_51_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg401_in = par_reset17_out ? 1'd0 : (right_52_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg401_write_en = (right_52_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_reset18_in = par_reset18_out ? 1'd0 : (par_done_reg402_out & par_done_reg403_out & par_done_reg404_out & par_done_reg405_out & par_done_reg406_out & par_done_reg407_out & par_done_reg408_out & par_done_reg409_out & par_done_reg410_out & par_done_reg411_out & par_done_reg412_out & par_done_reg413_out & par_done_reg414_out & par_done_reg415_out & par_done_reg416_out & par_done_reg417_out & par_done_reg418_out & par_done_reg419_out & par_done_reg420_out & par_done_reg421_out & par_done_reg422_out & par_done_reg423_out & par_done_reg424_out & par_done_reg425_out & par_done_reg426_out & par_done_reg427_out & par_done_reg428_out & par_done_reg429_out & par_done_reg430_out & par_done_reg431_out & par_done_reg432_out & par_done_reg433_out & par_done_reg434_out & par_done_reg435_out & par_done_reg436_out & par_done_reg437_out & par_done_reg438_out & par_done_reg439_out & par_done_reg440_out & par_done_reg441_out & par_done_reg442_out & par_done_reg443_out & par_done_reg444_out & par_done_reg445_out & par_done_reg446_out & par_done_reg447_out & par_done_reg448_out & par_done_reg449_out & par_done_reg450_out & par_done_reg451_out & par_done_reg452_out & par_done_reg453_out & par_done_reg454_out & par_done_reg455_out & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_reset18_write_en = (par_done_reg402_out & par_done_reg403_out & par_done_reg404_out & par_done_reg405_out & par_done_reg406_out & par_done_reg407_out & par_done_reg408_out & par_done_reg409_out & par_done_reg410_out & par_done_reg411_out & par_done_reg412_out & par_done_reg413_out & par_done_reg414_out & par_done_reg415_out & par_done_reg416_out & par_done_reg417_out & par_done_reg418_out & par_done_reg419_out & par_done_reg420_out & par_done_reg421_out & par_done_reg422_out & par_done_reg423_out & par_done_reg424_out & par_done_reg425_out & par_done_reg426_out & par_done_reg427_out & par_done_reg428_out & par_done_reg429_out & par_done_reg430_out & par_done_reg431_out & par_done_reg432_out & par_done_reg433_out & par_done_reg434_out & par_done_reg435_out & par_done_reg436_out & par_done_reg437_out & par_done_reg438_out & par_done_reg439_out & par_done_reg440_out & par_done_reg441_out & par_done_reg442_out & par_done_reg443_out & par_done_reg444_out & par_done_reg445_out & par_done_reg446_out & par_done_reg447_out & par_done_reg448_out & par_done_reg449_out & par_done_reg450_out & par_done_reg451_out & par_done_reg452_out & par_done_reg453_out & par_done_reg454_out & par_done_reg455_out & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg402_in = par_reset18_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg402_write_en = (top_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg403_in = par_reset18_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg403_write_en = (top_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg404_in = par_reset18_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg404_write_en = (top_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg405_in = par_reset18_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg405_write_en = (top_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg406_in = par_reset18_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg406_write_en = (top_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg407_in = par_reset18_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg407_write_en = (top_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg408_in = par_reset18_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg408_write_en = (top_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg409_in = par_reset18_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg409_write_en = (top_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg410_in = par_reset18_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg410_write_en = (top_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg411_in = par_reset18_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg411_write_en = (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg412_in = par_reset18_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg412_write_en = (top_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg413_in = par_reset18_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg413_write_en = (top_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg414_in = par_reset18_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg414_write_en = (top_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg415_in = par_reset18_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg415_write_en = (top_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg416_in = par_reset18_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg416_write_en = (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg417_in = par_reset18_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg417_write_en = (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg418_in = par_reset18_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg418_write_en = (top_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg419_in = par_reset18_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg419_write_en = (top_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg420_in = par_reset18_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg420_write_en = (top_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg421_in = par_reset18_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg421_write_en = (top_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg422_in = par_reset18_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg422_write_en = (top_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg423_in = par_reset18_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg423_write_en = (top_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg424_in = par_reset18_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg424_write_en = (top_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg425_in = par_reset18_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg425_write_en = (top_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg426_in = par_reset18_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg426_write_en = (top_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg427_in = par_reset18_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg427_write_en = (top_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg428_in = par_reset18_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg428_write_en = (top_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg429_in = par_reset18_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg429_write_en = (left_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg430_in = par_reset18_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg430_write_en = (left_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg431_in = par_reset18_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg431_write_en = (left_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg432_in = par_reset18_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg432_write_en = (left_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg433_in = par_reset18_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg433_write_en = (left_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg434_in = par_reset18_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg434_write_en = (left_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg435_in = par_reset18_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg435_write_en = (left_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg436_in = par_reset18_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg436_write_en = (left_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg437_in = par_reset18_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg437_write_en = (left_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg438_in = par_reset18_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg438_write_en = (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg439_in = par_reset18_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg439_write_en = (left_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg440_in = par_reset18_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg440_write_en = (left_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg441_in = par_reset18_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg441_write_en = (left_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg442_in = par_reset18_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg442_write_en = (left_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg443_in = par_reset18_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg443_write_en = (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg444_in = par_reset18_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg444_write_en = (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg445_in = par_reset18_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg445_write_en = (left_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg446_in = par_reset18_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg446_write_en = (left_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg447_in = par_reset18_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg447_write_en = (left_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg448_in = par_reset18_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg448_write_en = (left_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg449_in = par_reset18_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg449_write_en = (left_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg450_in = par_reset18_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg450_write_en = (left_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg451_in = par_reset18_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg451_write_en = (left_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg452_in = par_reset18_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg452_write_en = (left_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg453_in = par_reset18_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg453_write_en = (left_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg454_in = par_reset18_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg454_write_en = (left_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg455_in = par_reset18_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg455_write_en = (left_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_reset19_in = par_reset19_out ? 1'd0 : (par_done_reg456_out & par_done_reg457_out & par_done_reg458_out & par_done_reg459_out & par_done_reg460_out & par_done_reg461_out & par_done_reg462_out & par_done_reg463_out & par_done_reg464_out & par_done_reg465_out & par_done_reg466_out & par_done_reg467_out & par_done_reg468_out & par_done_reg469_out & par_done_reg470_out & par_done_reg471_out & par_done_reg472_out & par_done_reg473_out & par_done_reg474_out & par_done_reg475_out & par_done_reg476_out & par_done_reg477_out & par_done_reg478_out & par_done_reg479_out & par_done_reg480_out & par_done_reg481_out & par_done_reg482_out & par_done_reg483_out & par_done_reg484_out & par_done_reg485_out & par_done_reg486_out & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_reset19_write_en = (par_done_reg456_out & par_done_reg457_out & par_done_reg458_out & par_done_reg459_out & par_done_reg460_out & par_done_reg461_out & par_done_reg462_out & par_done_reg463_out & par_done_reg464_out & par_done_reg465_out & par_done_reg466_out & par_done_reg467_out & par_done_reg468_out & par_done_reg469_out & par_done_reg470_out & par_done_reg471_out & par_done_reg472_out & par_done_reg473_out & par_done_reg474_out & par_done_reg475_out & par_done_reg476_out & par_done_reg477_out & par_done_reg478_out & par_done_reg479_out & par_done_reg480_out & par_done_reg481_out & par_done_reg482_out & par_done_reg483_out & par_done_reg484_out & par_done_reg485_out & par_done_reg486_out & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg456_in = par_reset19_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg456_write_en = (t4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg457_in = par_reset19_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg457_write_en = (t5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg458_in = par_reset19_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg458_write_en = (l4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg459_in = par_reset19_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg459_write_en = (l5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg460_in = par_reset19_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg460_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg461_in = par_reset19_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg461_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg462_in = par_reset19_out ? 1'd0 : (down_05_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg462_write_en = (down_05_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg463_in = par_reset19_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg463_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg464_in = par_reset19_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg464_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg465_in = par_reset19_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg465_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg466_in = par_reset19_out ? 1'd0 : (down_15_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg466_write_en = (down_15_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg467_in = par_reset19_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg467_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg468_in = par_reset19_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg468_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg469_in = par_reset19_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg469_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg470_in = par_reset19_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg470_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg471_in = par_reset19_out ? 1'd0 : (down_25_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg471_write_en = (down_25_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg472_in = par_reset19_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg472_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg473_in = par_reset19_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg473_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg474_in = par_reset19_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg474_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg475_in = par_reset19_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg475_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg476_in = par_reset19_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg476_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg477_in = par_reset19_out ? 1'd0 : (down_35_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg477_write_en = (down_35_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg478_in = par_reset19_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg478_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg479_in = par_reset19_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg479_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg480_in = par_reset19_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg480_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg481_in = par_reset19_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg481_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg482_in = par_reset19_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg482_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg483_in = par_reset19_out ? 1'd0 : (right_50_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg483_write_en = (right_50_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg484_in = par_reset19_out ? 1'd0 : (right_51_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg484_write_en = (right_51_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg485_in = par_reset19_out ? 1'd0 : (right_52_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg485_write_en = (right_52_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg486_in = par_reset19_out ? 1'd0 : (right_53_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg486_write_en = (right_53_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_reset20_in = par_reset20_out ? 1'd0 : (par_done_reg487_out & par_done_reg488_out & par_done_reg489_out & par_done_reg490_out & par_done_reg491_out & par_done_reg492_out & par_done_reg493_out & par_done_reg494_out & par_done_reg495_out & par_done_reg496_out & par_done_reg497_out & par_done_reg498_out & par_done_reg499_out & par_done_reg500_out & par_done_reg501_out & par_done_reg502_out & par_done_reg503_out & par_done_reg504_out & par_done_reg505_out & par_done_reg506_out & par_done_reg507_out & par_done_reg508_out & par_done_reg509_out & par_done_reg510_out & par_done_reg511_out & par_done_reg512_out & par_done_reg513_out & par_done_reg514_out & par_done_reg515_out & par_done_reg516_out & par_done_reg517_out & par_done_reg518_out & par_done_reg519_out & par_done_reg520_out & par_done_reg521_out & par_done_reg522_out & par_done_reg523_out & par_done_reg524_out & par_done_reg525_out & par_done_reg526_out & par_done_reg527_out & par_done_reg528_out & par_done_reg529_out & par_done_reg530_out & par_done_reg531_out & par_done_reg532_out & par_done_reg533_out & par_done_reg534_out & par_done_reg535_out & par_done_reg536_out & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_reset20_write_en = (par_done_reg487_out & par_done_reg488_out & par_done_reg489_out & par_done_reg490_out & par_done_reg491_out & par_done_reg492_out & par_done_reg493_out & par_done_reg494_out & par_done_reg495_out & par_done_reg496_out & par_done_reg497_out & par_done_reg498_out & par_done_reg499_out & par_done_reg500_out & par_done_reg501_out & par_done_reg502_out & par_done_reg503_out & par_done_reg504_out & par_done_reg505_out & par_done_reg506_out & par_done_reg507_out & par_done_reg508_out & par_done_reg509_out & par_done_reg510_out & par_done_reg511_out & par_done_reg512_out & par_done_reg513_out & par_done_reg514_out & par_done_reg515_out & par_done_reg516_out & par_done_reg517_out & par_done_reg518_out & par_done_reg519_out & par_done_reg520_out & par_done_reg521_out & par_done_reg522_out & par_done_reg523_out & par_done_reg524_out & par_done_reg525_out & par_done_reg526_out & par_done_reg527_out & par_done_reg528_out & par_done_reg529_out & par_done_reg530_out & par_done_reg531_out & par_done_reg532_out & par_done_reg533_out & par_done_reg534_out & par_done_reg535_out & par_done_reg536_out & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg487_in = par_reset20_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg487_write_en = (top_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg488_in = par_reset20_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg488_write_en = (top_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg489_in = par_reset20_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg489_write_en = (top_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg490_in = par_reset20_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg490_write_en = (top_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg491_in = par_reset20_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg491_write_en = (top_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg492_in = par_reset20_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg492_write_en = (top_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg493_in = par_reset20_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg493_write_en = (top_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg494_in = par_reset20_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg494_write_en = (top_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg495_in = par_reset20_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg495_write_en = (top_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg496_in = par_reset20_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg496_write_en = (top_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg497_in = par_reset20_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg497_write_en = (top_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg498_in = par_reset20_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg498_write_en = (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg499_in = par_reset20_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg499_write_en = (top_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg500_in = par_reset20_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg500_write_en = (top_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg501_in = par_reset20_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg501_write_en = (top_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg502_in = par_reset20_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg502_write_en = (top_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg503_in = par_reset20_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg503_write_en = (top_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg504_in = par_reset20_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg504_write_en = (top_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg505_in = par_reset20_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg505_write_en = (top_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg506_in = par_reset20_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg506_write_en = (top_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg507_in = par_reset20_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg507_write_en = (top_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg508_in = par_reset20_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg508_write_en = (top_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg509_in = par_reset20_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg509_write_en = (top_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg510_in = par_reset20_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg510_write_en = (top_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg511_in = par_reset20_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg511_write_en = (top_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg512_in = par_reset20_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg512_write_en = (left_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg513_in = par_reset20_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg513_write_en = (left_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg514_in = par_reset20_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg514_write_en = (left_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg515_in = par_reset20_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg515_write_en = (left_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg516_in = par_reset20_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg516_write_en = (left_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg517_in = par_reset20_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg517_write_en = (left_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg518_in = par_reset20_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg518_write_en = (left_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg519_in = par_reset20_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg519_write_en = (left_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg520_in = par_reset20_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg520_write_en = (left_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg521_in = par_reset20_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg521_write_en = (left_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg522_in = par_reset20_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg522_write_en = (left_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg523_in = par_reset20_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg523_write_en = (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg524_in = par_reset20_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg524_write_en = (left_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg525_in = par_reset20_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg525_write_en = (left_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg526_in = par_reset20_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg526_write_en = (left_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg527_in = par_reset20_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg527_write_en = (left_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg528_in = par_reset20_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg528_write_en = (left_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg529_in = par_reset20_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg529_write_en = (left_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg530_in = par_reset20_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg530_write_en = (left_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg531_in = par_reset20_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg531_write_en = (left_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg532_in = par_reset20_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg532_write_en = (left_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg533_in = par_reset20_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg533_write_en = (left_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg534_in = par_reset20_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg534_write_en = (left_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg535_in = par_reset20_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg535_write_en = (left_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg536_in = par_reset20_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg536_write_en = (left_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_reset21_in = par_reset21_out ? 1'd0 : (par_done_reg537_out & par_done_reg538_out & par_done_reg539_out & par_done_reg540_out & par_done_reg541_out & par_done_reg542_out & par_done_reg543_out & par_done_reg544_out & par_done_reg545_out & par_done_reg546_out & par_done_reg547_out & par_done_reg548_out & par_done_reg549_out & par_done_reg550_out & par_done_reg551_out & par_done_reg552_out & par_done_reg553_out & par_done_reg554_out & par_done_reg555_out & par_done_reg556_out & par_done_reg557_out & par_done_reg558_out & par_done_reg559_out & par_done_reg560_out & par_done_reg561_out & par_done_reg562_out & par_done_reg563_out & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_reset21_write_en = (par_done_reg537_out & par_done_reg538_out & par_done_reg539_out & par_done_reg540_out & par_done_reg541_out & par_done_reg542_out & par_done_reg543_out & par_done_reg544_out & par_done_reg545_out & par_done_reg546_out & par_done_reg547_out & par_done_reg548_out & par_done_reg549_out & par_done_reg550_out & par_done_reg551_out & par_done_reg552_out & par_done_reg553_out & par_done_reg554_out & par_done_reg555_out & par_done_reg556_out & par_done_reg557_out & par_done_reg558_out & par_done_reg559_out & par_done_reg560_out & par_done_reg561_out & par_done_reg562_out & par_done_reg563_out & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg537_in = par_reset21_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg537_write_en = (t5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg538_in = par_reset21_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg538_write_en = (l5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg539_in = par_reset21_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg539_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg540_in = par_reset21_out ? 1'd0 : (down_05_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg540_write_en = (down_05_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg541_in = par_reset21_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg541_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg542_in = par_reset21_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg542_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg543_in = par_reset21_out ? 1'd0 : (down_15_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg543_write_en = (down_15_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg544_in = par_reset21_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg544_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg545_in = par_reset21_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg545_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg546_in = par_reset21_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg546_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg547_in = par_reset21_out ? 1'd0 : (down_25_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg547_write_en = (down_25_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg548_in = par_reset21_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg548_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg549_in = par_reset21_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg549_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg550_in = par_reset21_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg550_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg551_in = par_reset21_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg551_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg552_in = par_reset21_out ? 1'd0 : (down_35_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg552_write_en = (down_35_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg553_in = par_reset21_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg553_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg554_in = par_reset21_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg554_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg555_in = par_reset21_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg555_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg556_in = par_reset21_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg556_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg557_in = par_reset21_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg557_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg558_in = par_reset21_out ? 1'd0 : (down_45_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg558_write_en = (down_45_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg559_in = par_reset21_out ? 1'd0 : (right_50_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg559_write_en = (right_50_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg560_in = par_reset21_out ? 1'd0 : (right_51_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg560_write_en = (right_51_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg561_in = par_reset21_out ? 1'd0 : (right_52_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg561_write_en = (right_52_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg562_in = par_reset21_out ? 1'd0 : (right_53_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg562_write_en = (right_53_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg563_in = par_reset21_out ? 1'd0 : (right_54_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg563_write_en = (right_54_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_reset22_in = par_reset22_out ? 1'd0 : (par_done_reg564_out & par_done_reg565_out & par_done_reg566_out & par_done_reg567_out & par_done_reg568_out & par_done_reg569_out & par_done_reg570_out & par_done_reg571_out & par_done_reg572_out & par_done_reg573_out & par_done_reg574_out & par_done_reg575_out & par_done_reg576_out & par_done_reg577_out & par_done_reg578_out & par_done_reg579_out & par_done_reg580_out & par_done_reg581_out & par_done_reg582_out & par_done_reg583_out & par_done_reg584_out & par_done_reg585_out & par_done_reg586_out & par_done_reg587_out & par_done_reg588_out & par_done_reg589_out & par_done_reg590_out & par_done_reg591_out & par_done_reg592_out & par_done_reg593_out & par_done_reg594_out & par_done_reg595_out & par_done_reg596_out & par_done_reg597_out & par_done_reg598_out & par_done_reg599_out & par_done_reg600_out & par_done_reg601_out & par_done_reg602_out & par_done_reg603_out & par_done_reg604_out & par_done_reg605_out & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_reset22_write_en = (par_done_reg564_out & par_done_reg565_out & par_done_reg566_out & par_done_reg567_out & par_done_reg568_out & par_done_reg569_out & par_done_reg570_out & par_done_reg571_out & par_done_reg572_out & par_done_reg573_out & par_done_reg574_out & par_done_reg575_out & par_done_reg576_out & par_done_reg577_out & par_done_reg578_out & par_done_reg579_out & par_done_reg580_out & par_done_reg581_out & par_done_reg582_out & par_done_reg583_out & par_done_reg584_out & par_done_reg585_out & par_done_reg586_out & par_done_reg587_out & par_done_reg588_out & par_done_reg589_out & par_done_reg590_out & par_done_reg591_out & par_done_reg592_out & par_done_reg593_out & par_done_reg594_out & par_done_reg595_out & par_done_reg596_out & par_done_reg597_out & par_done_reg598_out & par_done_reg599_out & par_done_reg600_out & par_done_reg601_out & par_done_reg602_out & par_done_reg603_out & par_done_reg604_out & par_done_reg605_out & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg564_in = par_reset22_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg564_write_en = (top_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg565_in = par_reset22_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg565_write_en = (top_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg566_in = par_reset22_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg566_write_en = (top_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg567_in = par_reset22_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg567_write_en = (top_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg568_in = par_reset22_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg568_write_en = (top_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg569_in = par_reset22_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg569_write_en = (top_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg570_in = par_reset22_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg570_write_en = (top_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg571_in = par_reset22_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg571_write_en = (top_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg572_in = par_reset22_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg572_write_en = (top_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg573_in = par_reset22_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg573_write_en = (top_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg574_in = par_reset22_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg574_write_en = (top_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg575_in = par_reset22_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg575_write_en = (top_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg576_in = par_reset22_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg576_write_en = (top_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg577_in = par_reset22_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg577_write_en = (top_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg578_in = par_reset22_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg578_write_en = (top_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg579_in = par_reset22_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg579_write_en = (top_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg580_in = par_reset22_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg580_write_en = (top_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg581_in = par_reset22_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg581_write_en = (top_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg582_in = par_reset22_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg582_write_en = (top_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg583_in = par_reset22_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg583_write_en = (top_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg584_in = par_reset22_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg584_write_en = (top_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg585_in = par_reset22_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg585_write_en = (left_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg586_in = par_reset22_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg586_write_en = (left_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg587_in = par_reset22_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg587_write_en = (left_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg588_in = par_reset22_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg588_write_en = (left_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg589_in = par_reset22_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg589_write_en = (left_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg590_in = par_reset22_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg590_write_en = (left_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg591_in = par_reset22_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg591_write_en = (left_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg592_in = par_reset22_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg592_write_en = (left_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg593_in = par_reset22_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg593_write_en = (left_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg594_in = par_reset22_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg594_write_en = (left_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg595_in = par_reset22_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg595_write_en = (left_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg596_in = par_reset22_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg596_write_en = (left_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg597_in = par_reset22_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg597_write_en = (left_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg598_in = par_reset22_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg598_write_en = (left_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg599_in = par_reset22_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg599_write_en = (left_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg600_in = par_reset22_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg600_write_en = (left_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg601_in = par_reset22_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg601_write_en = (left_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg602_in = par_reset22_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg602_write_en = (left_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg603_in = par_reset22_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg603_write_en = (left_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg604_in = par_reset22_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg604_write_en = (left_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg605_in = par_reset22_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg605_write_en = (left_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_reset23_in = par_reset23_out ? 1'd0 : (par_done_reg606_out & par_done_reg607_out & par_done_reg608_out & par_done_reg609_out & par_done_reg610_out & par_done_reg611_out & par_done_reg612_out & par_done_reg613_out & par_done_reg614_out & par_done_reg615_out & par_done_reg616_out & par_done_reg617_out & par_done_reg618_out & par_done_reg619_out & par_done_reg620_out & par_done_reg621_out & par_done_reg622_out & par_done_reg623_out & par_done_reg624_out & par_done_reg625_out & par_done_reg626_out & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_reset23_write_en = (par_done_reg606_out & par_done_reg607_out & par_done_reg608_out & par_done_reg609_out & par_done_reg610_out & par_done_reg611_out & par_done_reg612_out & par_done_reg613_out & par_done_reg614_out & par_done_reg615_out & par_done_reg616_out & par_done_reg617_out & par_done_reg618_out & par_done_reg619_out & par_done_reg620_out & par_done_reg621_out & par_done_reg622_out & par_done_reg623_out & par_done_reg624_out & par_done_reg625_out & par_done_reg626_out & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg606_in = par_reset23_out ? 1'd0 : (down_05_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg606_write_en = (down_05_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg607_in = par_reset23_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg607_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg608_in = par_reset23_out ? 1'd0 : (down_15_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg608_write_en = (down_15_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg609_in = par_reset23_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg609_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg610_in = par_reset23_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg610_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg611_in = par_reset23_out ? 1'd0 : (down_25_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg611_write_en = (down_25_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg612_in = par_reset23_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg612_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg613_in = par_reset23_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg613_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg614_in = par_reset23_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg614_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg615_in = par_reset23_out ? 1'd0 : (down_35_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg615_write_en = (down_35_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg616_in = par_reset23_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg616_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg617_in = par_reset23_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg617_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg618_in = par_reset23_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg618_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg619_in = par_reset23_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg619_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg620_in = par_reset23_out ? 1'd0 : (down_45_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg620_write_en = (down_45_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg621_in = par_reset23_out ? 1'd0 : (right_50_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg621_write_en = (right_50_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg622_in = par_reset23_out ? 1'd0 : (right_51_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg622_write_en = (right_51_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg623_in = par_reset23_out ? 1'd0 : (right_52_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg623_write_en = (right_52_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg624_in = par_reset23_out ? 1'd0 : (right_53_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg624_write_en = (right_53_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg625_in = par_reset23_out ? 1'd0 : (right_54_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg625_write_en = (right_54_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg626_in = par_reset23_out ? 1'd0 : (pe_55_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg626_write_en = (pe_55_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_reset24_in = par_reset24_out ? 1'd0 : (par_done_reg627_out & par_done_reg628_out & par_done_reg629_out & par_done_reg630_out & par_done_reg631_out & par_done_reg632_out & par_done_reg633_out & par_done_reg634_out & par_done_reg635_out & par_done_reg636_out & par_done_reg637_out & par_done_reg638_out & par_done_reg639_out & par_done_reg640_out & par_done_reg641_out & par_done_reg642_out & par_done_reg643_out & par_done_reg644_out & par_done_reg645_out & par_done_reg646_out & par_done_reg647_out & par_done_reg648_out & par_done_reg649_out & par_done_reg650_out & par_done_reg651_out & par_done_reg652_out & par_done_reg653_out & par_done_reg654_out & par_done_reg655_out & par_done_reg656_out & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_reset24_write_en = (par_done_reg627_out & par_done_reg628_out & par_done_reg629_out & par_done_reg630_out & par_done_reg631_out & par_done_reg632_out & par_done_reg633_out & par_done_reg634_out & par_done_reg635_out & par_done_reg636_out & par_done_reg637_out & par_done_reg638_out & par_done_reg639_out & par_done_reg640_out & par_done_reg641_out & par_done_reg642_out & par_done_reg643_out & par_done_reg644_out & par_done_reg645_out & par_done_reg646_out & par_done_reg647_out & par_done_reg648_out & par_done_reg649_out & par_done_reg650_out & par_done_reg651_out & par_done_reg652_out & par_done_reg653_out & par_done_reg654_out & par_done_reg655_out & par_done_reg656_out & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg627_in = par_reset24_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg627_write_en = (top_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg628_in = par_reset24_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg628_write_en = (top_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg629_in = par_reset24_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg629_write_en = (top_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg630_in = par_reset24_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg630_write_en = (top_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg631_in = par_reset24_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg631_write_en = (top_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg632_in = par_reset24_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg632_write_en = (top_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg633_in = par_reset24_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg633_write_en = (top_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg634_in = par_reset24_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg634_write_en = (top_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg635_in = par_reset24_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg635_write_en = (top_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg636_in = par_reset24_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg636_write_en = (top_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg637_in = par_reset24_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg637_write_en = (top_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg638_in = par_reset24_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg638_write_en = (top_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg639_in = par_reset24_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg639_write_en = (top_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg640_in = par_reset24_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg640_write_en = (top_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg641_in = par_reset24_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg641_write_en = (top_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg642_in = par_reset24_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg642_write_en = (left_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg643_in = par_reset24_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg643_write_en = (left_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg644_in = par_reset24_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg644_write_en = (left_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg645_in = par_reset24_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg645_write_en = (left_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg646_in = par_reset24_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg646_write_en = (left_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg647_in = par_reset24_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg647_write_en = (left_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg648_in = par_reset24_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg648_write_en = (left_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg649_in = par_reset24_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg649_write_en = (left_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg650_in = par_reset24_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg650_write_en = (left_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg651_in = par_reset24_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg651_write_en = (left_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg652_in = par_reset24_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg652_write_en = (left_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg653_in = par_reset24_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg653_write_en = (left_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg654_in = par_reset24_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg654_write_en = (left_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg655_in = par_reset24_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg655_write_en = (left_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg656_in = par_reset24_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg656_write_en = (left_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_reset25_in = par_reset25_out ? 1'd0 : (par_done_reg657_out & par_done_reg658_out & par_done_reg659_out & par_done_reg660_out & par_done_reg661_out & par_done_reg662_out & par_done_reg663_out & par_done_reg664_out & par_done_reg665_out & par_done_reg666_out & par_done_reg667_out & par_done_reg668_out & par_done_reg669_out & par_done_reg670_out & par_done_reg671_out & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_reset25_write_en = (par_done_reg657_out & par_done_reg658_out & par_done_reg659_out & par_done_reg660_out & par_done_reg661_out & par_done_reg662_out & par_done_reg663_out & par_done_reg664_out & par_done_reg665_out & par_done_reg666_out & par_done_reg667_out & par_done_reg668_out & par_done_reg669_out & par_done_reg670_out & par_done_reg671_out & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg657_in = par_reset25_out ? 1'd0 : (down_15_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg657_write_en = (down_15_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg658_in = par_reset25_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg658_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg659_in = par_reset25_out ? 1'd0 : (down_25_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg659_write_en = (down_25_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg660_in = par_reset25_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg660_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg661_in = par_reset25_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg661_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg662_in = par_reset25_out ? 1'd0 : (down_35_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg662_write_en = (down_35_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg663_in = par_reset25_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg663_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg664_in = par_reset25_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg664_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg665_in = par_reset25_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg665_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg666_in = par_reset25_out ? 1'd0 : (down_45_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg666_write_en = (down_45_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg667_in = par_reset25_out ? 1'd0 : (right_51_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg667_write_en = (right_51_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg668_in = par_reset25_out ? 1'd0 : (right_52_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg668_write_en = (right_52_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg669_in = par_reset25_out ? 1'd0 : (right_53_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg669_write_en = (right_53_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg670_in = par_reset25_out ? 1'd0 : (right_54_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg670_write_en = (right_54_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg671_in = par_reset25_out ? 1'd0 : (pe_55_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg671_write_en = (pe_55_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_reset26_in = par_reset26_out ? 1'd0 : (par_done_reg672_out & par_done_reg673_out & par_done_reg674_out & par_done_reg675_out & par_done_reg676_out & par_done_reg677_out & par_done_reg678_out & par_done_reg679_out & par_done_reg680_out & par_done_reg681_out & par_done_reg682_out & par_done_reg683_out & par_done_reg684_out & par_done_reg685_out & par_done_reg686_out & par_done_reg687_out & par_done_reg688_out & par_done_reg689_out & par_done_reg690_out & par_done_reg691_out & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_reset26_write_en = (par_done_reg672_out & par_done_reg673_out & par_done_reg674_out & par_done_reg675_out & par_done_reg676_out & par_done_reg677_out & par_done_reg678_out & par_done_reg679_out & par_done_reg680_out & par_done_reg681_out & par_done_reg682_out & par_done_reg683_out & par_done_reg684_out & par_done_reg685_out & par_done_reg686_out & par_done_reg687_out & par_done_reg688_out & par_done_reg689_out & par_done_reg690_out & par_done_reg691_out & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg672_in = par_reset26_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg672_write_en = (top_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg673_in = par_reset26_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg673_write_en = (top_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg674_in = par_reset26_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg674_write_en = (top_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg675_in = par_reset26_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg675_write_en = (top_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg676_in = par_reset26_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg676_write_en = (top_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg677_in = par_reset26_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg677_write_en = (top_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg678_in = par_reset26_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg678_write_en = (top_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg679_in = par_reset26_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg679_write_en = (top_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg680_in = par_reset26_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg680_write_en = (top_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg681_in = par_reset26_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg681_write_en = (top_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg682_in = par_reset26_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg682_write_en = (left_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg683_in = par_reset26_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg683_write_en = (left_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg684_in = par_reset26_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg684_write_en = (left_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg685_in = par_reset26_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg685_write_en = (left_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg686_in = par_reset26_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg686_write_en = (left_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg687_in = par_reset26_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg687_write_en = (left_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg688_in = par_reset26_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg688_write_en = (left_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg689_in = par_reset26_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg689_write_en = (left_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg690_in = par_reset26_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg690_write_en = (left_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg691_in = par_reset26_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg691_write_en = (left_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_reset27_in = par_reset27_out ? 1'd0 : (par_done_reg692_out & par_done_reg693_out & par_done_reg694_out & par_done_reg695_out & par_done_reg696_out & par_done_reg697_out & par_done_reg698_out & par_done_reg699_out & par_done_reg700_out & par_done_reg701_out & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_reset27_write_en = (par_done_reg692_out & par_done_reg693_out & par_done_reg694_out & par_done_reg695_out & par_done_reg696_out & par_done_reg697_out & par_done_reg698_out & par_done_reg699_out & par_done_reg700_out & par_done_reg701_out & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg692_in = par_reset27_out ? 1'd0 : (down_25_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg692_write_en = (down_25_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg693_in = par_reset27_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg693_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg694_in = par_reset27_out ? 1'd0 : (down_35_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg694_write_en = (down_35_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg695_in = par_reset27_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg695_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg696_in = par_reset27_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg696_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg697_in = par_reset27_out ? 1'd0 : (down_45_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg697_write_en = (down_45_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg698_in = par_reset27_out ? 1'd0 : (right_52_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg698_write_en = (right_52_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg699_in = par_reset27_out ? 1'd0 : (right_53_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg699_write_en = (right_53_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg700_in = par_reset27_out ? 1'd0 : (right_54_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg700_write_en = (right_54_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg701_in = par_reset27_out ? 1'd0 : (pe_55_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg701_write_en = (pe_55_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_reset28_in = par_reset28_out ? 1'd0 : (par_done_reg702_out & par_done_reg703_out & par_done_reg704_out & par_done_reg705_out & par_done_reg706_out & par_done_reg707_out & par_done_reg708_out & par_done_reg709_out & par_done_reg710_out & par_done_reg711_out & par_done_reg712_out & par_done_reg713_out & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_reset28_write_en = (par_done_reg702_out & par_done_reg703_out & par_done_reg704_out & par_done_reg705_out & par_done_reg706_out & par_done_reg707_out & par_done_reg708_out & par_done_reg709_out & par_done_reg710_out & par_done_reg711_out & par_done_reg712_out & par_done_reg713_out & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg702_in = par_reset28_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg702_write_en = (top_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg703_in = par_reset28_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg703_write_en = (top_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg704_in = par_reset28_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg704_write_en = (top_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg705_in = par_reset28_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg705_write_en = (top_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg706_in = par_reset28_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg706_write_en = (top_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg707_in = par_reset28_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg707_write_en = (top_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg708_in = par_reset28_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg708_write_en = (left_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg709_in = par_reset28_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg709_write_en = (left_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg710_in = par_reset28_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg710_write_en = (left_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg711_in = par_reset28_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg711_write_en = (left_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg712_in = par_reset28_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg712_write_en = (left_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg713_in = par_reset28_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg713_write_en = (left_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_reset29_in = par_reset29_out ? 1'd0 : (par_done_reg714_out & par_done_reg715_out & par_done_reg716_out & par_done_reg717_out & par_done_reg718_out & par_done_reg719_out & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_reset29_write_en = (par_done_reg714_out & par_done_reg715_out & par_done_reg716_out & par_done_reg717_out & par_done_reg718_out & par_done_reg719_out & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg714_in = par_reset29_out ? 1'd0 : (down_35_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg714_write_en = (down_35_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg715_in = par_reset29_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg715_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg716_in = par_reset29_out ? 1'd0 : (down_45_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg716_write_en = (down_45_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg717_in = par_reset29_out ? 1'd0 : (right_53_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg717_write_en = (right_53_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg718_in = par_reset29_out ? 1'd0 : (right_54_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg718_write_en = (right_54_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg719_in = par_reset29_out ? 1'd0 : (pe_55_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg719_write_en = (pe_55_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_reset30_in = par_reset30_out ? 1'd0 : (par_done_reg720_out & par_done_reg721_out & par_done_reg722_out & par_done_reg723_out & par_done_reg724_out & par_done_reg725_out & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_reset30_write_en = (par_done_reg720_out & par_done_reg721_out & par_done_reg722_out & par_done_reg723_out & par_done_reg724_out & par_done_reg725_out & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg720_in = par_reset30_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg720_write_en = (top_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg721_in = par_reset30_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg721_write_en = (top_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg722_in = par_reset30_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg722_write_en = (top_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg723_in = par_reset30_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg723_write_en = (left_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg724_in = par_reset30_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg724_write_en = (left_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg725_in = par_reset30_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg725_write_en = (left_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_reset31_in = par_reset31_out ? 1'd0 : (par_done_reg726_out & par_done_reg727_out & par_done_reg728_out & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_reset31_write_en = (par_done_reg726_out & par_done_reg727_out & par_done_reg728_out & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg726_in = par_reset31_out ? 1'd0 : (down_45_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg726_write_en = (down_45_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg727_in = par_reset31_out ? 1'd0 : (right_54_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg727_write_en = (right_54_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg728_in = par_reset31_out ? 1'd0 : (pe_55_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg728_write_en = (pe_55_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_reset32_in = par_reset32_out ? 1'd0 : (par_done_reg729_out & par_done_reg730_out & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_reset32_write_en = (par_done_reg729_out & par_done_reg730_out & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg729_in = par_reset32_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg729_write_en = (top_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg730_in = par_reset32_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg730_write_en = (left_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_reset33_in = par_reset33_out ? 1'd0 : (par_done_reg731_out & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_reset33_write_en = (par_done_reg731_out & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg731_in = par_reset33_out ? 1'd0 : (pe_55_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg731_write_en = (pe_55_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd70) ? 32'd0 : (fsm0_out == 32'd69 & out_mem_done & go) ? 32'd70 : (fsm0_out == 32'd68 & out_mem_done & go) ? 32'd69 : (fsm0_out == 32'd67 & out_mem_done & go) ? 32'd68 : (fsm0_out == 32'd66 & out_mem_done & go) ? 32'd67 : (fsm0_out == 32'd65 & out_mem_done & go) ? 32'd66 : (fsm0_out == 32'd64 & out_mem_done & go) ? 32'd65 : (fsm0_out == 32'd63 & out_mem_done & go) ? 32'd64 : (fsm0_out == 32'd62 & out_mem_done & go) ? 32'd63 : (fsm0_out == 32'd61 & out_mem_done & go) ? 32'd62 : (fsm0_out == 32'd60 & out_mem_done & go) ? 32'd61 : (fsm0_out == 32'd59 & out_mem_done & go) ? 32'd60 : (fsm0_out == 32'd58 & out_mem_done & go) ? 32'd59 : (fsm0_out == 32'd57 & out_mem_done & go) ? 32'd58 : (fsm0_out == 32'd56 & out_mem_done & go) ? 32'd57 : (fsm0_out == 32'd55 & out_mem_done & go) ? 32'd56 : (fsm0_out == 32'd54 & out_mem_done & go) ? 32'd55 : (fsm0_out == 32'd53 & out_mem_done & go) ? 32'd54 : (fsm0_out == 32'd52 & out_mem_done & go) ? 32'd53 : (fsm0_out == 32'd51 & out_mem_done & go) ? 32'd52 : (fsm0_out == 32'd50 & out_mem_done & go) ? 32'd51 : (fsm0_out == 32'd49 & out_mem_done & go) ? 32'd50 : (fsm0_out == 32'd48 & out_mem_done & go) ? 32'd49 : (fsm0_out == 32'd47 & out_mem_done & go) ? 32'd48 : (fsm0_out == 32'd46 & out_mem_done & go) ? 32'd47 : (fsm0_out == 32'd45 & out_mem_done & go) ? 32'd46 : (fsm0_out == 32'd44 & out_mem_done & go) ? 32'd45 : (fsm0_out == 32'd43 & out_mem_done & go) ? 32'd44 : (fsm0_out == 32'd42 & out_mem_done & go) ? 32'd43 : (fsm0_out == 32'd41 & out_mem_done & go) ? 32'd42 : (fsm0_out == 32'd40 & out_mem_done & go) ? 32'd41 : (fsm0_out == 32'd39 & out_mem_done & go) ? 32'd40 : (fsm0_out == 32'd38 & out_mem_done & go) ? 32'd39 : (fsm0_out == 32'd37 & out_mem_done & go) ? 32'd38 : (fsm0_out == 32'd36 & out_mem_done & go) ? 32'd37 : (fsm0_out == 32'd35 & out_mem_done & go) ? 32'd36 : (fsm0_out == 32'd34 & out_mem_done & go) ? 32'd35 : (fsm0_out == 32'd33 & par_reset33_out & go) ? 32'd34 : (fsm0_out == 32'd32 & par_reset32_out & go) ? 32'd33 : (fsm0_out == 32'd31 & par_reset31_out & go) ? 32'd32 : (fsm0_out == 32'd30 & par_reset30_out & go) ? 32'd31 : (fsm0_out == 32'd29 & par_reset29_out & go) ? 32'd30 : (fsm0_out == 32'd28 & par_reset28_out & go) ? 32'd29 : (fsm0_out == 32'd27 & par_reset27_out & go) ? 32'd28 : (fsm0_out == 32'd26 & par_reset26_out & go) ? 32'd27 : (fsm0_out == 32'd25 & par_reset25_out & go) ? 32'd26 : (fsm0_out == 32'd24 & par_reset24_out & go) ? 32'd25 : (fsm0_out == 32'd23 & par_reset23_out & go) ? 32'd24 : (fsm0_out == 32'd22 & par_reset22_out & go) ? 32'd23 : (fsm0_out == 32'd21 & par_reset21_out & go) ? 32'd22 : (fsm0_out == 32'd20 & par_reset20_out & go) ? 32'd21 : (fsm0_out == 32'd19 & par_reset19_out & go) ? 32'd20 : (fsm0_out == 32'd18 & par_reset18_out & go) ? 32'd19 : (fsm0_out == 32'd17 & par_reset17_out & go) ? 32'd18 : (fsm0_out == 32'd16 & par_reset16_out & go) ? 32'd17 : (fsm0_out == 32'd15 & par_reset15_out & go) ? 32'd16 : (fsm0_out == 32'd14 & par_reset14_out & go) ? 32'd15 : (fsm0_out == 32'd13 & par_reset13_out & go) ? 32'd14 : (fsm0_out == 32'd12 & par_reset12_out & go) ? 32'd13 : (fsm0_out == 32'd11 & par_reset11_out & go) ? 32'd12 : (fsm0_out == 32'd10 & par_reset10_out & go) ? 32'd11 : (fsm0_out == 32'd9 & par_reset9_out & go) ? 32'd10 : (fsm0_out == 32'd8 & par_reset8_out & go) ? 32'd9 : (fsm0_out == 32'd7 & par_reset7_out & go) ? 32'd8 : (fsm0_out == 32'd6 & par_reset6_out & go) ? 32'd7 : (fsm0_out == 32'd5 & par_reset5_out & go) ? 32'd6 : (fsm0_out == 32'd4 & par_reset4_out & go) ? 32'd5 : (fsm0_out == 32'd3 & par_reset3_out & go) ? 32'd4 : (fsm0_out == 32'd2 & par_reset2_out & go) ? 32'd3 : (fsm0_out == 32'd1 & par_reset1_out & go) ? 32'd2 : (fsm0_out == 32'd0 & par_reset0_out & go) ? 32'd1 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & par_reset0_out & go | fsm0_out == 32'd1 & par_reset1_out & go | fsm0_out == 32'd2 & par_reset2_out & go | fsm0_out == 32'd3 & par_reset3_out & go | fsm0_out == 32'd4 & par_reset4_out & go | fsm0_out == 32'd5 & par_reset5_out & go | fsm0_out == 32'd6 & par_reset6_out & go | fsm0_out == 32'd7 & par_reset7_out & go | fsm0_out == 32'd8 & par_reset8_out & go | fsm0_out == 32'd9 & par_reset9_out & go | fsm0_out == 32'd10 & par_reset10_out & go | fsm0_out == 32'd11 & par_reset11_out & go | fsm0_out == 32'd12 & par_reset12_out & go | fsm0_out == 32'd13 & par_reset13_out & go | fsm0_out == 32'd14 & par_reset14_out & go | fsm0_out == 32'd15 & par_reset15_out & go | fsm0_out == 32'd16 & par_reset16_out & go | fsm0_out == 32'd17 & par_reset17_out & go | fsm0_out == 32'd18 & par_reset18_out & go | fsm0_out == 32'd19 & par_reset19_out & go | fsm0_out == 32'd20 & par_reset20_out & go | fsm0_out == 32'd21 & par_reset21_out & go | fsm0_out == 32'd22 & par_reset22_out & go | fsm0_out == 32'd23 & par_reset23_out & go | fsm0_out == 32'd24 & par_reset24_out & go | fsm0_out == 32'd25 & par_reset25_out & go | fsm0_out == 32'd26 & par_reset26_out & go | fsm0_out == 32'd27 & par_reset27_out & go | fsm0_out == 32'd28 & par_reset28_out & go | fsm0_out == 32'd29 & par_reset29_out & go | fsm0_out == 32'd30 & par_reset30_out & go | fsm0_out == 32'd31 & par_reset31_out & go | fsm0_out == 32'd32 & par_reset32_out & go | fsm0_out == 32'd33 & par_reset33_out & go | fsm0_out == 32'd34 & out_mem_done & go | fsm0_out == 32'd35 & out_mem_done & go | fsm0_out == 32'd36 & out_mem_done & go | fsm0_out == 32'd37 & out_mem_done & go | fsm0_out == 32'd38 & out_mem_done & go | fsm0_out == 32'd39 & out_mem_done & go | fsm0_out == 32'd40 & out_mem_done & go | fsm0_out == 32'd41 & out_mem_done & go | fsm0_out == 32'd42 & out_mem_done & go | fsm0_out == 32'd43 & out_mem_done & go | fsm0_out == 32'd44 & out_mem_done & go | fsm0_out == 32'd45 & out_mem_done & go | fsm0_out == 32'd46 & out_mem_done & go | fsm0_out == 32'd47 & out_mem_done & go | fsm0_out == 32'd48 & out_mem_done & go | fsm0_out == 32'd49 & out_mem_done & go | fsm0_out == 32'd50 & out_mem_done & go | fsm0_out == 32'd51 & out_mem_done & go | fsm0_out == 32'd52 & out_mem_done & go | fsm0_out == 32'd53 & out_mem_done & go | fsm0_out == 32'd54 & out_mem_done & go | fsm0_out == 32'd55 & out_mem_done & go | fsm0_out == 32'd56 & out_mem_done & go | fsm0_out == 32'd57 & out_mem_done & go | fsm0_out == 32'd58 & out_mem_done & go | fsm0_out == 32'd59 & out_mem_done & go | fsm0_out == 32'd60 & out_mem_done & go | fsm0_out == 32'd61 & out_mem_done & go | fsm0_out == 32'd62 & out_mem_done & go | fsm0_out == 32'd63 & out_mem_done & go | fsm0_out == 32'd64 & out_mem_done & go | fsm0_out == 32'd65 & out_mem_done & go | fsm0_out == 32'd66 & out_mem_done & go | fsm0_out == 32'd67 & out_mem_done & go | fsm0_out == 32'd68 & out_mem_done & go | fsm0_out == 32'd69 & out_mem_done & go | fsm0_out == 32'd70) ? 1'd1 : '0;
endmodule // end main