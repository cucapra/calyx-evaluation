/* verilator lint_off WIDTH */
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule

module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule

module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule

// Component Signature
module mac_pe (
      input wire [31:0] top,
      input wire [31:0] left,
      input wire go,
      input wire clk,
      output wire [31:0] down,
      output wire [31:0] right,
      output wire [31:0] out,
      output wire done
  );
  
  // Structure wire declarations
  wire [31:0] mul_left;
  wire [31:0] mul_right;
  wire mul_go;
  wire mul_clk;
  wire [31:0] mul_out;
  wire mul_done;
  wire [31:0] add_left;
  wire [31:0] add_right;
  wire [31:0] add_out;
  wire [31:0] mul_reg_in;
  wire mul_reg_write_en;
  wire mul_reg_clk;
  wire [31:0] mul_reg_out;
  wire mul_reg_done;
  wire [31:0] acc_in;
  wire acc_write_en;
  wire acc_clk;
  wire [31:0] acc_out;
  wire acc_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_mult_pipe #(32) mul (
      .left(mul_left),
      .right(mul_right),
      .go(mul_go),
      .clk(clk),
      .out(mul_out),
      .done(mul_done)
  );
  
  std_add #(32) add (
      .left(add_left),
      .right(add_right),
      .out(add_out)
  );
  
  std_reg #(32) mul_reg (
      .in(mul_reg_in),
      .write_en(mul_reg_write_en),
      .clk(clk),
      .out(mul_reg_out),
      .done(mul_reg_done)
  );
  
  std_reg #(32) acc (
      .in(acc_in),
      .write_en(acc_write_en),
      .clk(clk),
      .out(acc_out),
      .done(acc_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign down = top;
  assign right = left;
  assign out = acc_out;
  assign done = (fsm0_out == 32'd2) ? 1'd1 : '0;
  assign mul_left = (fsm0_out == 32'd0 & !mul_reg_done & go) ? top : '0;
  assign mul_right = (fsm0_out == 32'd0 & !mul_reg_done & go) ? left : '0;
  assign mul_go = (!mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign add_left = (fsm0_out == 32'd1 & !acc_done & go) ? acc_out : '0;
  assign add_right = (fsm0_out == 32'd1 & !acc_done & go) ? mul_reg_out : '0;
  assign mul_reg_in = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? mul_out : '0;
  assign mul_reg_write_en = (mul_done & fsm0_out == 32'd0 & !mul_reg_done & go) ? 1'd1 : '0;
  assign acc_in = (fsm0_out == 32'd1 & !acc_done & go) ? add_out : '0;
  assign acc_write_en = (fsm0_out == 32'd1 & !acc_done & go) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd1 & acc_done & go) ? 32'd2 : (fsm0_out == 32'd0 & mul_reg_done & go) ? 32'd1 : (fsm0_out == 32'd2) ? 32'd0 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & mul_reg_done & go | fsm0_out == 32'd1 & acc_done & go | fsm0_out == 32'd2) ? 1'd1 : '0;
endmodule // end mac_pe
// Component Signature
module main (
      input wire go,
      input wire clk,
      input wire [31:0] out_mem_read_data,
      input wire out_mem_done,
      output wire done,
      output wire [3:0] out_mem_addr0,
      output wire [3:0] out_mem_addr1,
      output wire [31:0] out_mem_write_data,
      output wire out_mem_write_en
  );
  
  // Structure wire declarations
  wire [31:0] left_77_read_in;
  wire left_77_read_write_en;
  wire left_77_read_clk;
  wire [31:0] left_77_read_out;
  wire left_77_read_done;
  wire [31:0] top_77_read_in;
  wire top_77_read_write_en;
  wire top_77_read_clk;
  wire [31:0] top_77_read_out;
  wire top_77_read_done;
  wire [31:0] pe_77_top;
  wire [31:0] pe_77_left;
  wire pe_77_go;
  wire pe_77_clk;
  wire [31:0] pe_77_down;
  wire [31:0] pe_77_right;
  wire [31:0] pe_77_out;
  wire pe_77_done;
  wire [31:0] right_76_write_in;
  wire right_76_write_write_en;
  wire right_76_write_clk;
  wire [31:0] right_76_write_out;
  wire right_76_write_done;
  wire [31:0] left_76_read_in;
  wire left_76_read_write_en;
  wire left_76_read_clk;
  wire [31:0] left_76_read_out;
  wire left_76_read_done;
  wire [31:0] top_76_read_in;
  wire top_76_read_write_en;
  wire top_76_read_clk;
  wire [31:0] top_76_read_out;
  wire top_76_read_done;
  wire [31:0] pe_76_top;
  wire [31:0] pe_76_left;
  wire pe_76_go;
  wire pe_76_clk;
  wire [31:0] pe_76_down;
  wire [31:0] pe_76_right;
  wire [31:0] pe_76_out;
  wire pe_76_done;
  wire [31:0] right_75_write_in;
  wire right_75_write_write_en;
  wire right_75_write_clk;
  wire [31:0] right_75_write_out;
  wire right_75_write_done;
  wire [31:0] left_75_read_in;
  wire left_75_read_write_en;
  wire left_75_read_clk;
  wire [31:0] left_75_read_out;
  wire left_75_read_done;
  wire [31:0] top_75_read_in;
  wire top_75_read_write_en;
  wire top_75_read_clk;
  wire [31:0] top_75_read_out;
  wire top_75_read_done;
  wire [31:0] pe_75_top;
  wire [31:0] pe_75_left;
  wire pe_75_go;
  wire pe_75_clk;
  wire [31:0] pe_75_down;
  wire [31:0] pe_75_right;
  wire [31:0] pe_75_out;
  wire pe_75_done;
  wire [31:0] right_74_write_in;
  wire right_74_write_write_en;
  wire right_74_write_clk;
  wire [31:0] right_74_write_out;
  wire right_74_write_done;
  wire [31:0] left_74_read_in;
  wire left_74_read_write_en;
  wire left_74_read_clk;
  wire [31:0] left_74_read_out;
  wire left_74_read_done;
  wire [31:0] top_74_read_in;
  wire top_74_read_write_en;
  wire top_74_read_clk;
  wire [31:0] top_74_read_out;
  wire top_74_read_done;
  wire [31:0] pe_74_top;
  wire [31:0] pe_74_left;
  wire pe_74_go;
  wire pe_74_clk;
  wire [31:0] pe_74_down;
  wire [31:0] pe_74_right;
  wire [31:0] pe_74_out;
  wire pe_74_done;
  wire [31:0] right_73_write_in;
  wire right_73_write_write_en;
  wire right_73_write_clk;
  wire [31:0] right_73_write_out;
  wire right_73_write_done;
  wire [31:0] left_73_read_in;
  wire left_73_read_write_en;
  wire left_73_read_clk;
  wire [31:0] left_73_read_out;
  wire left_73_read_done;
  wire [31:0] top_73_read_in;
  wire top_73_read_write_en;
  wire top_73_read_clk;
  wire [31:0] top_73_read_out;
  wire top_73_read_done;
  wire [31:0] pe_73_top;
  wire [31:0] pe_73_left;
  wire pe_73_go;
  wire pe_73_clk;
  wire [31:0] pe_73_down;
  wire [31:0] pe_73_right;
  wire [31:0] pe_73_out;
  wire pe_73_done;
  wire [31:0] right_72_write_in;
  wire right_72_write_write_en;
  wire right_72_write_clk;
  wire [31:0] right_72_write_out;
  wire right_72_write_done;
  wire [31:0] left_72_read_in;
  wire left_72_read_write_en;
  wire left_72_read_clk;
  wire [31:0] left_72_read_out;
  wire left_72_read_done;
  wire [31:0] top_72_read_in;
  wire top_72_read_write_en;
  wire top_72_read_clk;
  wire [31:0] top_72_read_out;
  wire top_72_read_done;
  wire [31:0] pe_72_top;
  wire [31:0] pe_72_left;
  wire pe_72_go;
  wire pe_72_clk;
  wire [31:0] pe_72_down;
  wire [31:0] pe_72_right;
  wire [31:0] pe_72_out;
  wire pe_72_done;
  wire [31:0] right_71_write_in;
  wire right_71_write_write_en;
  wire right_71_write_clk;
  wire [31:0] right_71_write_out;
  wire right_71_write_done;
  wire [31:0] left_71_read_in;
  wire left_71_read_write_en;
  wire left_71_read_clk;
  wire [31:0] left_71_read_out;
  wire left_71_read_done;
  wire [31:0] top_71_read_in;
  wire top_71_read_write_en;
  wire top_71_read_clk;
  wire [31:0] top_71_read_out;
  wire top_71_read_done;
  wire [31:0] pe_71_top;
  wire [31:0] pe_71_left;
  wire pe_71_go;
  wire pe_71_clk;
  wire [31:0] pe_71_down;
  wire [31:0] pe_71_right;
  wire [31:0] pe_71_out;
  wire pe_71_done;
  wire [31:0] right_70_write_in;
  wire right_70_write_write_en;
  wire right_70_write_clk;
  wire [31:0] right_70_write_out;
  wire right_70_write_done;
  wire [31:0] left_70_read_in;
  wire left_70_read_write_en;
  wire left_70_read_clk;
  wire [31:0] left_70_read_out;
  wire left_70_read_done;
  wire [31:0] top_70_read_in;
  wire top_70_read_write_en;
  wire top_70_read_clk;
  wire [31:0] top_70_read_out;
  wire top_70_read_done;
  wire [31:0] pe_70_top;
  wire [31:0] pe_70_left;
  wire pe_70_go;
  wire pe_70_clk;
  wire [31:0] pe_70_down;
  wire [31:0] pe_70_right;
  wire [31:0] pe_70_out;
  wire pe_70_done;
  wire [31:0] down_67_write_in;
  wire down_67_write_write_en;
  wire down_67_write_clk;
  wire [31:0] down_67_write_out;
  wire down_67_write_done;
  wire [31:0] left_67_read_in;
  wire left_67_read_write_en;
  wire left_67_read_clk;
  wire [31:0] left_67_read_out;
  wire left_67_read_done;
  wire [31:0] top_67_read_in;
  wire top_67_read_write_en;
  wire top_67_read_clk;
  wire [31:0] top_67_read_out;
  wire top_67_read_done;
  wire [31:0] pe_67_top;
  wire [31:0] pe_67_left;
  wire pe_67_go;
  wire pe_67_clk;
  wire [31:0] pe_67_down;
  wire [31:0] pe_67_right;
  wire [31:0] pe_67_out;
  wire pe_67_done;
  wire [31:0] down_66_write_in;
  wire down_66_write_write_en;
  wire down_66_write_clk;
  wire [31:0] down_66_write_out;
  wire down_66_write_done;
  wire [31:0] right_66_write_in;
  wire right_66_write_write_en;
  wire right_66_write_clk;
  wire [31:0] right_66_write_out;
  wire right_66_write_done;
  wire [31:0] left_66_read_in;
  wire left_66_read_write_en;
  wire left_66_read_clk;
  wire [31:0] left_66_read_out;
  wire left_66_read_done;
  wire [31:0] top_66_read_in;
  wire top_66_read_write_en;
  wire top_66_read_clk;
  wire [31:0] top_66_read_out;
  wire top_66_read_done;
  wire [31:0] pe_66_top;
  wire [31:0] pe_66_left;
  wire pe_66_go;
  wire pe_66_clk;
  wire [31:0] pe_66_down;
  wire [31:0] pe_66_right;
  wire [31:0] pe_66_out;
  wire pe_66_done;
  wire [31:0] down_65_write_in;
  wire down_65_write_write_en;
  wire down_65_write_clk;
  wire [31:0] down_65_write_out;
  wire down_65_write_done;
  wire [31:0] right_65_write_in;
  wire right_65_write_write_en;
  wire right_65_write_clk;
  wire [31:0] right_65_write_out;
  wire right_65_write_done;
  wire [31:0] left_65_read_in;
  wire left_65_read_write_en;
  wire left_65_read_clk;
  wire [31:0] left_65_read_out;
  wire left_65_read_done;
  wire [31:0] top_65_read_in;
  wire top_65_read_write_en;
  wire top_65_read_clk;
  wire [31:0] top_65_read_out;
  wire top_65_read_done;
  wire [31:0] pe_65_top;
  wire [31:0] pe_65_left;
  wire pe_65_go;
  wire pe_65_clk;
  wire [31:0] pe_65_down;
  wire [31:0] pe_65_right;
  wire [31:0] pe_65_out;
  wire pe_65_done;
  wire [31:0] down_64_write_in;
  wire down_64_write_write_en;
  wire down_64_write_clk;
  wire [31:0] down_64_write_out;
  wire down_64_write_done;
  wire [31:0] right_64_write_in;
  wire right_64_write_write_en;
  wire right_64_write_clk;
  wire [31:0] right_64_write_out;
  wire right_64_write_done;
  wire [31:0] left_64_read_in;
  wire left_64_read_write_en;
  wire left_64_read_clk;
  wire [31:0] left_64_read_out;
  wire left_64_read_done;
  wire [31:0] top_64_read_in;
  wire top_64_read_write_en;
  wire top_64_read_clk;
  wire [31:0] top_64_read_out;
  wire top_64_read_done;
  wire [31:0] pe_64_top;
  wire [31:0] pe_64_left;
  wire pe_64_go;
  wire pe_64_clk;
  wire [31:0] pe_64_down;
  wire [31:0] pe_64_right;
  wire [31:0] pe_64_out;
  wire pe_64_done;
  wire [31:0] down_63_write_in;
  wire down_63_write_write_en;
  wire down_63_write_clk;
  wire [31:0] down_63_write_out;
  wire down_63_write_done;
  wire [31:0] right_63_write_in;
  wire right_63_write_write_en;
  wire right_63_write_clk;
  wire [31:0] right_63_write_out;
  wire right_63_write_done;
  wire [31:0] left_63_read_in;
  wire left_63_read_write_en;
  wire left_63_read_clk;
  wire [31:0] left_63_read_out;
  wire left_63_read_done;
  wire [31:0] top_63_read_in;
  wire top_63_read_write_en;
  wire top_63_read_clk;
  wire [31:0] top_63_read_out;
  wire top_63_read_done;
  wire [31:0] pe_63_top;
  wire [31:0] pe_63_left;
  wire pe_63_go;
  wire pe_63_clk;
  wire [31:0] pe_63_down;
  wire [31:0] pe_63_right;
  wire [31:0] pe_63_out;
  wire pe_63_done;
  wire [31:0] down_62_write_in;
  wire down_62_write_write_en;
  wire down_62_write_clk;
  wire [31:0] down_62_write_out;
  wire down_62_write_done;
  wire [31:0] right_62_write_in;
  wire right_62_write_write_en;
  wire right_62_write_clk;
  wire [31:0] right_62_write_out;
  wire right_62_write_done;
  wire [31:0] left_62_read_in;
  wire left_62_read_write_en;
  wire left_62_read_clk;
  wire [31:0] left_62_read_out;
  wire left_62_read_done;
  wire [31:0] top_62_read_in;
  wire top_62_read_write_en;
  wire top_62_read_clk;
  wire [31:0] top_62_read_out;
  wire top_62_read_done;
  wire [31:0] pe_62_top;
  wire [31:0] pe_62_left;
  wire pe_62_go;
  wire pe_62_clk;
  wire [31:0] pe_62_down;
  wire [31:0] pe_62_right;
  wire [31:0] pe_62_out;
  wire pe_62_done;
  wire [31:0] down_61_write_in;
  wire down_61_write_write_en;
  wire down_61_write_clk;
  wire [31:0] down_61_write_out;
  wire down_61_write_done;
  wire [31:0] right_61_write_in;
  wire right_61_write_write_en;
  wire right_61_write_clk;
  wire [31:0] right_61_write_out;
  wire right_61_write_done;
  wire [31:0] left_61_read_in;
  wire left_61_read_write_en;
  wire left_61_read_clk;
  wire [31:0] left_61_read_out;
  wire left_61_read_done;
  wire [31:0] top_61_read_in;
  wire top_61_read_write_en;
  wire top_61_read_clk;
  wire [31:0] top_61_read_out;
  wire top_61_read_done;
  wire [31:0] pe_61_top;
  wire [31:0] pe_61_left;
  wire pe_61_go;
  wire pe_61_clk;
  wire [31:0] pe_61_down;
  wire [31:0] pe_61_right;
  wire [31:0] pe_61_out;
  wire pe_61_done;
  wire [31:0] down_60_write_in;
  wire down_60_write_write_en;
  wire down_60_write_clk;
  wire [31:0] down_60_write_out;
  wire down_60_write_done;
  wire [31:0] right_60_write_in;
  wire right_60_write_write_en;
  wire right_60_write_clk;
  wire [31:0] right_60_write_out;
  wire right_60_write_done;
  wire [31:0] left_60_read_in;
  wire left_60_read_write_en;
  wire left_60_read_clk;
  wire [31:0] left_60_read_out;
  wire left_60_read_done;
  wire [31:0] top_60_read_in;
  wire top_60_read_write_en;
  wire top_60_read_clk;
  wire [31:0] top_60_read_out;
  wire top_60_read_done;
  wire [31:0] pe_60_top;
  wire [31:0] pe_60_left;
  wire pe_60_go;
  wire pe_60_clk;
  wire [31:0] pe_60_down;
  wire [31:0] pe_60_right;
  wire [31:0] pe_60_out;
  wire pe_60_done;
  wire [31:0] down_57_write_in;
  wire down_57_write_write_en;
  wire down_57_write_clk;
  wire [31:0] down_57_write_out;
  wire down_57_write_done;
  wire [31:0] left_57_read_in;
  wire left_57_read_write_en;
  wire left_57_read_clk;
  wire [31:0] left_57_read_out;
  wire left_57_read_done;
  wire [31:0] top_57_read_in;
  wire top_57_read_write_en;
  wire top_57_read_clk;
  wire [31:0] top_57_read_out;
  wire top_57_read_done;
  wire [31:0] pe_57_top;
  wire [31:0] pe_57_left;
  wire pe_57_go;
  wire pe_57_clk;
  wire [31:0] pe_57_down;
  wire [31:0] pe_57_right;
  wire [31:0] pe_57_out;
  wire pe_57_done;
  wire [31:0] down_56_write_in;
  wire down_56_write_write_en;
  wire down_56_write_clk;
  wire [31:0] down_56_write_out;
  wire down_56_write_done;
  wire [31:0] right_56_write_in;
  wire right_56_write_write_en;
  wire right_56_write_clk;
  wire [31:0] right_56_write_out;
  wire right_56_write_done;
  wire [31:0] left_56_read_in;
  wire left_56_read_write_en;
  wire left_56_read_clk;
  wire [31:0] left_56_read_out;
  wire left_56_read_done;
  wire [31:0] top_56_read_in;
  wire top_56_read_write_en;
  wire top_56_read_clk;
  wire [31:0] top_56_read_out;
  wire top_56_read_done;
  wire [31:0] pe_56_top;
  wire [31:0] pe_56_left;
  wire pe_56_go;
  wire pe_56_clk;
  wire [31:0] pe_56_down;
  wire [31:0] pe_56_right;
  wire [31:0] pe_56_out;
  wire pe_56_done;
  wire [31:0] down_55_write_in;
  wire down_55_write_write_en;
  wire down_55_write_clk;
  wire [31:0] down_55_write_out;
  wire down_55_write_done;
  wire [31:0] right_55_write_in;
  wire right_55_write_write_en;
  wire right_55_write_clk;
  wire [31:0] right_55_write_out;
  wire right_55_write_done;
  wire [31:0] left_55_read_in;
  wire left_55_read_write_en;
  wire left_55_read_clk;
  wire [31:0] left_55_read_out;
  wire left_55_read_done;
  wire [31:0] top_55_read_in;
  wire top_55_read_write_en;
  wire top_55_read_clk;
  wire [31:0] top_55_read_out;
  wire top_55_read_done;
  wire [31:0] pe_55_top;
  wire [31:0] pe_55_left;
  wire pe_55_go;
  wire pe_55_clk;
  wire [31:0] pe_55_down;
  wire [31:0] pe_55_right;
  wire [31:0] pe_55_out;
  wire pe_55_done;
  wire [31:0] down_54_write_in;
  wire down_54_write_write_en;
  wire down_54_write_clk;
  wire [31:0] down_54_write_out;
  wire down_54_write_done;
  wire [31:0] right_54_write_in;
  wire right_54_write_write_en;
  wire right_54_write_clk;
  wire [31:0] right_54_write_out;
  wire right_54_write_done;
  wire [31:0] left_54_read_in;
  wire left_54_read_write_en;
  wire left_54_read_clk;
  wire [31:0] left_54_read_out;
  wire left_54_read_done;
  wire [31:0] top_54_read_in;
  wire top_54_read_write_en;
  wire top_54_read_clk;
  wire [31:0] top_54_read_out;
  wire top_54_read_done;
  wire [31:0] pe_54_top;
  wire [31:0] pe_54_left;
  wire pe_54_go;
  wire pe_54_clk;
  wire [31:0] pe_54_down;
  wire [31:0] pe_54_right;
  wire [31:0] pe_54_out;
  wire pe_54_done;
  wire [31:0] down_53_write_in;
  wire down_53_write_write_en;
  wire down_53_write_clk;
  wire [31:0] down_53_write_out;
  wire down_53_write_done;
  wire [31:0] right_53_write_in;
  wire right_53_write_write_en;
  wire right_53_write_clk;
  wire [31:0] right_53_write_out;
  wire right_53_write_done;
  wire [31:0] left_53_read_in;
  wire left_53_read_write_en;
  wire left_53_read_clk;
  wire [31:0] left_53_read_out;
  wire left_53_read_done;
  wire [31:0] top_53_read_in;
  wire top_53_read_write_en;
  wire top_53_read_clk;
  wire [31:0] top_53_read_out;
  wire top_53_read_done;
  wire [31:0] pe_53_top;
  wire [31:0] pe_53_left;
  wire pe_53_go;
  wire pe_53_clk;
  wire [31:0] pe_53_down;
  wire [31:0] pe_53_right;
  wire [31:0] pe_53_out;
  wire pe_53_done;
  wire [31:0] down_52_write_in;
  wire down_52_write_write_en;
  wire down_52_write_clk;
  wire [31:0] down_52_write_out;
  wire down_52_write_done;
  wire [31:0] right_52_write_in;
  wire right_52_write_write_en;
  wire right_52_write_clk;
  wire [31:0] right_52_write_out;
  wire right_52_write_done;
  wire [31:0] left_52_read_in;
  wire left_52_read_write_en;
  wire left_52_read_clk;
  wire [31:0] left_52_read_out;
  wire left_52_read_done;
  wire [31:0] top_52_read_in;
  wire top_52_read_write_en;
  wire top_52_read_clk;
  wire [31:0] top_52_read_out;
  wire top_52_read_done;
  wire [31:0] pe_52_top;
  wire [31:0] pe_52_left;
  wire pe_52_go;
  wire pe_52_clk;
  wire [31:0] pe_52_down;
  wire [31:0] pe_52_right;
  wire [31:0] pe_52_out;
  wire pe_52_done;
  wire [31:0] down_51_write_in;
  wire down_51_write_write_en;
  wire down_51_write_clk;
  wire [31:0] down_51_write_out;
  wire down_51_write_done;
  wire [31:0] right_51_write_in;
  wire right_51_write_write_en;
  wire right_51_write_clk;
  wire [31:0] right_51_write_out;
  wire right_51_write_done;
  wire [31:0] left_51_read_in;
  wire left_51_read_write_en;
  wire left_51_read_clk;
  wire [31:0] left_51_read_out;
  wire left_51_read_done;
  wire [31:0] top_51_read_in;
  wire top_51_read_write_en;
  wire top_51_read_clk;
  wire [31:0] top_51_read_out;
  wire top_51_read_done;
  wire [31:0] pe_51_top;
  wire [31:0] pe_51_left;
  wire pe_51_go;
  wire pe_51_clk;
  wire [31:0] pe_51_down;
  wire [31:0] pe_51_right;
  wire [31:0] pe_51_out;
  wire pe_51_done;
  wire [31:0] down_50_write_in;
  wire down_50_write_write_en;
  wire down_50_write_clk;
  wire [31:0] down_50_write_out;
  wire down_50_write_done;
  wire [31:0] right_50_write_in;
  wire right_50_write_write_en;
  wire right_50_write_clk;
  wire [31:0] right_50_write_out;
  wire right_50_write_done;
  wire [31:0] left_50_read_in;
  wire left_50_read_write_en;
  wire left_50_read_clk;
  wire [31:0] left_50_read_out;
  wire left_50_read_done;
  wire [31:0] top_50_read_in;
  wire top_50_read_write_en;
  wire top_50_read_clk;
  wire [31:0] top_50_read_out;
  wire top_50_read_done;
  wire [31:0] pe_50_top;
  wire [31:0] pe_50_left;
  wire pe_50_go;
  wire pe_50_clk;
  wire [31:0] pe_50_down;
  wire [31:0] pe_50_right;
  wire [31:0] pe_50_out;
  wire pe_50_done;
  wire [31:0] down_47_write_in;
  wire down_47_write_write_en;
  wire down_47_write_clk;
  wire [31:0] down_47_write_out;
  wire down_47_write_done;
  wire [31:0] left_47_read_in;
  wire left_47_read_write_en;
  wire left_47_read_clk;
  wire [31:0] left_47_read_out;
  wire left_47_read_done;
  wire [31:0] top_47_read_in;
  wire top_47_read_write_en;
  wire top_47_read_clk;
  wire [31:0] top_47_read_out;
  wire top_47_read_done;
  wire [31:0] pe_47_top;
  wire [31:0] pe_47_left;
  wire pe_47_go;
  wire pe_47_clk;
  wire [31:0] pe_47_down;
  wire [31:0] pe_47_right;
  wire [31:0] pe_47_out;
  wire pe_47_done;
  wire [31:0] down_46_write_in;
  wire down_46_write_write_en;
  wire down_46_write_clk;
  wire [31:0] down_46_write_out;
  wire down_46_write_done;
  wire [31:0] right_46_write_in;
  wire right_46_write_write_en;
  wire right_46_write_clk;
  wire [31:0] right_46_write_out;
  wire right_46_write_done;
  wire [31:0] left_46_read_in;
  wire left_46_read_write_en;
  wire left_46_read_clk;
  wire [31:0] left_46_read_out;
  wire left_46_read_done;
  wire [31:0] top_46_read_in;
  wire top_46_read_write_en;
  wire top_46_read_clk;
  wire [31:0] top_46_read_out;
  wire top_46_read_done;
  wire [31:0] pe_46_top;
  wire [31:0] pe_46_left;
  wire pe_46_go;
  wire pe_46_clk;
  wire [31:0] pe_46_down;
  wire [31:0] pe_46_right;
  wire [31:0] pe_46_out;
  wire pe_46_done;
  wire [31:0] down_45_write_in;
  wire down_45_write_write_en;
  wire down_45_write_clk;
  wire [31:0] down_45_write_out;
  wire down_45_write_done;
  wire [31:0] right_45_write_in;
  wire right_45_write_write_en;
  wire right_45_write_clk;
  wire [31:0] right_45_write_out;
  wire right_45_write_done;
  wire [31:0] left_45_read_in;
  wire left_45_read_write_en;
  wire left_45_read_clk;
  wire [31:0] left_45_read_out;
  wire left_45_read_done;
  wire [31:0] top_45_read_in;
  wire top_45_read_write_en;
  wire top_45_read_clk;
  wire [31:0] top_45_read_out;
  wire top_45_read_done;
  wire [31:0] pe_45_top;
  wire [31:0] pe_45_left;
  wire pe_45_go;
  wire pe_45_clk;
  wire [31:0] pe_45_down;
  wire [31:0] pe_45_right;
  wire [31:0] pe_45_out;
  wire pe_45_done;
  wire [31:0] down_44_write_in;
  wire down_44_write_write_en;
  wire down_44_write_clk;
  wire [31:0] down_44_write_out;
  wire down_44_write_done;
  wire [31:0] right_44_write_in;
  wire right_44_write_write_en;
  wire right_44_write_clk;
  wire [31:0] right_44_write_out;
  wire right_44_write_done;
  wire [31:0] left_44_read_in;
  wire left_44_read_write_en;
  wire left_44_read_clk;
  wire [31:0] left_44_read_out;
  wire left_44_read_done;
  wire [31:0] top_44_read_in;
  wire top_44_read_write_en;
  wire top_44_read_clk;
  wire [31:0] top_44_read_out;
  wire top_44_read_done;
  wire [31:0] pe_44_top;
  wire [31:0] pe_44_left;
  wire pe_44_go;
  wire pe_44_clk;
  wire [31:0] pe_44_down;
  wire [31:0] pe_44_right;
  wire [31:0] pe_44_out;
  wire pe_44_done;
  wire [31:0] down_43_write_in;
  wire down_43_write_write_en;
  wire down_43_write_clk;
  wire [31:0] down_43_write_out;
  wire down_43_write_done;
  wire [31:0] right_43_write_in;
  wire right_43_write_write_en;
  wire right_43_write_clk;
  wire [31:0] right_43_write_out;
  wire right_43_write_done;
  wire [31:0] left_43_read_in;
  wire left_43_read_write_en;
  wire left_43_read_clk;
  wire [31:0] left_43_read_out;
  wire left_43_read_done;
  wire [31:0] top_43_read_in;
  wire top_43_read_write_en;
  wire top_43_read_clk;
  wire [31:0] top_43_read_out;
  wire top_43_read_done;
  wire [31:0] pe_43_top;
  wire [31:0] pe_43_left;
  wire pe_43_go;
  wire pe_43_clk;
  wire [31:0] pe_43_down;
  wire [31:0] pe_43_right;
  wire [31:0] pe_43_out;
  wire pe_43_done;
  wire [31:0] down_42_write_in;
  wire down_42_write_write_en;
  wire down_42_write_clk;
  wire [31:0] down_42_write_out;
  wire down_42_write_done;
  wire [31:0] right_42_write_in;
  wire right_42_write_write_en;
  wire right_42_write_clk;
  wire [31:0] right_42_write_out;
  wire right_42_write_done;
  wire [31:0] left_42_read_in;
  wire left_42_read_write_en;
  wire left_42_read_clk;
  wire [31:0] left_42_read_out;
  wire left_42_read_done;
  wire [31:0] top_42_read_in;
  wire top_42_read_write_en;
  wire top_42_read_clk;
  wire [31:0] top_42_read_out;
  wire top_42_read_done;
  wire [31:0] pe_42_top;
  wire [31:0] pe_42_left;
  wire pe_42_go;
  wire pe_42_clk;
  wire [31:0] pe_42_down;
  wire [31:0] pe_42_right;
  wire [31:0] pe_42_out;
  wire pe_42_done;
  wire [31:0] down_41_write_in;
  wire down_41_write_write_en;
  wire down_41_write_clk;
  wire [31:0] down_41_write_out;
  wire down_41_write_done;
  wire [31:0] right_41_write_in;
  wire right_41_write_write_en;
  wire right_41_write_clk;
  wire [31:0] right_41_write_out;
  wire right_41_write_done;
  wire [31:0] left_41_read_in;
  wire left_41_read_write_en;
  wire left_41_read_clk;
  wire [31:0] left_41_read_out;
  wire left_41_read_done;
  wire [31:0] top_41_read_in;
  wire top_41_read_write_en;
  wire top_41_read_clk;
  wire [31:0] top_41_read_out;
  wire top_41_read_done;
  wire [31:0] pe_41_top;
  wire [31:0] pe_41_left;
  wire pe_41_go;
  wire pe_41_clk;
  wire [31:0] pe_41_down;
  wire [31:0] pe_41_right;
  wire [31:0] pe_41_out;
  wire pe_41_done;
  wire [31:0] down_40_write_in;
  wire down_40_write_write_en;
  wire down_40_write_clk;
  wire [31:0] down_40_write_out;
  wire down_40_write_done;
  wire [31:0] right_40_write_in;
  wire right_40_write_write_en;
  wire right_40_write_clk;
  wire [31:0] right_40_write_out;
  wire right_40_write_done;
  wire [31:0] left_40_read_in;
  wire left_40_read_write_en;
  wire left_40_read_clk;
  wire [31:0] left_40_read_out;
  wire left_40_read_done;
  wire [31:0] top_40_read_in;
  wire top_40_read_write_en;
  wire top_40_read_clk;
  wire [31:0] top_40_read_out;
  wire top_40_read_done;
  wire [31:0] pe_40_top;
  wire [31:0] pe_40_left;
  wire pe_40_go;
  wire pe_40_clk;
  wire [31:0] pe_40_down;
  wire [31:0] pe_40_right;
  wire [31:0] pe_40_out;
  wire pe_40_done;
  wire [31:0] down_37_write_in;
  wire down_37_write_write_en;
  wire down_37_write_clk;
  wire [31:0] down_37_write_out;
  wire down_37_write_done;
  wire [31:0] left_37_read_in;
  wire left_37_read_write_en;
  wire left_37_read_clk;
  wire [31:0] left_37_read_out;
  wire left_37_read_done;
  wire [31:0] top_37_read_in;
  wire top_37_read_write_en;
  wire top_37_read_clk;
  wire [31:0] top_37_read_out;
  wire top_37_read_done;
  wire [31:0] pe_37_top;
  wire [31:0] pe_37_left;
  wire pe_37_go;
  wire pe_37_clk;
  wire [31:0] pe_37_down;
  wire [31:0] pe_37_right;
  wire [31:0] pe_37_out;
  wire pe_37_done;
  wire [31:0] down_36_write_in;
  wire down_36_write_write_en;
  wire down_36_write_clk;
  wire [31:0] down_36_write_out;
  wire down_36_write_done;
  wire [31:0] right_36_write_in;
  wire right_36_write_write_en;
  wire right_36_write_clk;
  wire [31:0] right_36_write_out;
  wire right_36_write_done;
  wire [31:0] left_36_read_in;
  wire left_36_read_write_en;
  wire left_36_read_clk;
  wire [31:0] left_36_read_out;
  wire left_36_read_done;
  wire [31:0] top_36_read_in;
  wire top_36_read_write_en;
  wire top_36_read_clk;
  wire [31:0] top_36_read_out;
  wire top_36_read_done;
  wire [31:0] pe_36_top;
  wire [31:0] pe_36_left;
  wire pe_36_go;
  wire pe_36_clk;
  wire [31:0] pe_36_down;
  wire [31:0] pe_36_right;
  wire [31:0] pe_36_out;
  wire pe_36_done;
  wire [31:0] down_35_write_in;
  wire down_35_write_write_en;
  wire down_35_write_clk;
  wire [31:0] down_35_write_out;
  wire down_35_write_done;
  wire [31:0] right_35_write_in;
  wire right_35_write_write_en;
  wire right_35_write_clk;
  wire [31:0] right_35_write_out;
  wire right_35_write_done;
  wire [31:0] left_35_read_in;
  wire left_35_read_write_en;
  wire left_35_read_clk;
  wire [31:0] left_35_read_out;
  wire left_35_read_done;
  wire [31:0] top_35_read_in;
  wire top_35_read_write_en;
  wire top_35_read_clk;
  wire [31:0] top_35_read_out;
  wire top_35_read_done;
  wire [31:0] pe_35_top;
  wire [31:0] pe_35_left;
  wire pe_35_go;
  wire pe_35_clk;
  wire [31:0] pe_35_down;
  wire [31:0] pe_35_right;
  wire [31:0] pe_35_out;
  wire pe_35_done;
  wire [31:0] down_34_write_in;
  wire down_34_write_write_en;
  wire down_34_write_clk;
  wire [31:0] down_34_write_out;
  wire down_34_write_done;
  wire [31:0] right_34_write_in;
  wire right_34_write_write_en;
  wire right_34_write_clk;
  wire [31:0] right_34_write_out;
  wire right_34_write_done;
  wire [31:0] left_34_read_in;
  wire left_34_read_write_en;
  wire left_34_read_clk;
  wire [31:0] left_34_read_out;
  wire left_34_read_done;
  wire [31:0] top_34_read_in;
  wire top_34_read_write_en;
  wire top_34_read_clk;
  wire [31:0] top_34_read_out;
  wire top_34_read_done;
  wire [31:0] pe_34_top;
  wire [31:0] pe_34_left;
  wire pe_34_go;
  wire pe_34_clk;
  wire [31:0] pe_34_down;
  wire [31:0] pe_34_right;
  wire [31:0] pe_34_out;
  wire pe_34_done;
  wire [31:0] down_33_write_in;
  wire down_33_write_write_en;
  wire down_33_write_clk;
  wire [31:0] down_33_write_out;
  wire down_33_write_done;
  wire [31:0] right_33_write_in;
  wire right_33_write_write_en;
  wire right_33_write_clk;
  wire [31:0] right_33_write_out;
  wire right_33_write_done;
  wire [31:0] left_33_read_in;
  wire left_33_read_write_en;
  wire left_33_read_clk;
  wire [31:0] left_33_read_out;
  wire left_33_read_done;
  wire [31:0] top_33_read_in;
  wire top_33_read_write_en;
  wire top_33_read_clk;
  wire [31:0] top_33_read_out;
  wire top_33_read_done;
  wire [31:0] pe_33_top;
  wire [31:0] pe_33_left;
  wire pe_33_go;
  wire pe_33_clk;
  wire [31:0] pe_33_down;
  wire [31:0] pe_33_right;
  wire [31:0] pe_33_out;
  wire pe_33_done;
  wire [31:0] down_32_write_in;
  wire down_32_write_write_en;
  wire down_32_write_clk;
  wire [31:0] down_32_write_out;
  wire down_32_write_done;
  wire [31:0] right_32_write_in;
  wire right_32_write_write_en;
  wire right_32_write_clk;
  wire [31:0] right_32_write_out;
  wire right_32_write_done;
  wire [31:0] left_32_read_in;
  wire left_32_read_write_en;
  wire left_32_read_clk;
  wire [31:0] left_32_read_out;
  wire left_32_read_done;
  wire [31:0] top_32_read_in;
  wire top_32_read_write_en;
  wire top_32_read_clk;
  wire [31:0] top_32_read_out;
  wire top_32_read_done;
  wire [31:0] pe_32_top;
  wire [31:0] pe_32_left;
  wire pe_32_go;
  wire pe_32_clk;
  wire [31:0] pe_32_down;
  wire [31:0] pe_32_right;
  wire [31:0] pe_32_out;
  wire pe_32_done;
  wire [31:0] down_31_write_in;
  wire down_31_write_write_en;
  wire down_31_write_clk;
  wire [31:0] down_31_write_out;
  wire down_31_write_done;
  wire [31:0] right_31_write_in;
  wire right_31_write_write_en;
  wire right_31_write_clk;
  wire [31:0] right_31_write_out;
  wire right_31_write_done;
  wire [31:0] left_31_read_in;
  wire left_31_read_write_en;
  wire left_31_read_clk;
  wire [31:0] left_31_read_out;
  wire left_31_read_done;
  wire [31:0] top_31_read_in;
  wire top_31_read_write_en;
  wire top_31_read_clk;
  wire [31:0] top_31_read_out;
  wire top_31_read_done;
  wire [31:0] pe_31_top;
  wire [31:0] pe_31_left;
  wire pe_31_go;
  wire pe_31_clk;
  wire [31:0] pe_31_down;
  wire [31:0] pe_31_right;
  wire [31:0] pe_31_out;
  wire pe_31_done;
  wire [31:0] down_30_write_in;
  wire down_30_write_write_en;
  wire down_30_write_clk;
  wire [31:0] down_30_write_out;
  wire down_30_write_done;
  wire [31:0] right_30_write_in;
  wire right_30_write_write_en;
  wire right_30_write_clk;
  wire [31:0] right_30_write_out;
  wire right_30_write_done;
  wire [31:0] left_30_read_in;
  wire left_30_read_write_en;
  wire left_30_read_clk;
  wire [31:0] left_30_read_out;
  wire left_30_read_done;
  wire [31:0] top_30_read_in;
  wire top_30_read_write_en;
  wire top_30_read_clk;
  wire [31:0] top_30_read_out;
  wire top_30_read_done;
  wire [31:0] pe_30_top;
  wire [31:0] pe_30_left;
  wire pe_30_go;
  wire pe_30_clk;
  wire [31:0] pe_30_down;
  wire [31:0] pe_30_right;
  wire [31:0] pe_30_out;
  wire pe_30_done;
  wire [31:0] down_27_write_in;
  wire down_27_write_write_en;
  wire down_27_write_clk;
  wire [31:0] down_27_write_out;
  wire down_27_write_done;
  wire [31:0] left_27_read_in;
  wire left_27_read_write_en;
  wire left_27_read_clk;
  wire [31:0] left_27_read_out;
  wire left_27_read_done;
  wire [31:0] top_27_read_in;
  wire top_27_read_write_en;
  wire top_27_read_clk;
  wire [31:0] top_27_read_out;
  wire top_27_read_done;
  wire [31:0] pe_27_top;
  wire [31:0] pe_27_left;
  wire pe_27_go;
  wire pe_27_clk;
  wire [31:0] pe_27_down;
  wire [31:0] pe_27_right;
  wire [31:0] pe_27_out;
  wire pe_27_done;
  wire [31:0] down_26_write_in;
  wire down_26_write_write_en;
  wire down_26_write_clk;
  wire [31:0] down_26_write_out;
  wire down_26_write_done;
  wire [31:0] right_26_write_in;
  wire right_26_write_write_en;
  wire right_26_write_clk;
  wire [31:0] right_26_write_out;
  wire right_26_write_done;
  wire [31:0] left_26_read_in;
  wire left_26_read_write_en;
  wire left_26_read_clk;
  wire [31:0] left_26_read_out;
  wire left_26_read_done;
  wire [31:0] top_26_read_in;
  wire top_26_read_write_en;
  wire top_26_read_clk;
  wire [31:0] top_26_read_out;
  wire top_26_read_done;
  wire [31:0] pe_26_top;
  wire [31:0] pe_26_left;
  wire pe_26_go;
  wire pe_26_clk;
  wire [31:0] pe_26_down;
  wire [31:0] pe_26_right;
  wire [31:0] pe_26_out;
  wire pe_26_done;
  wire [31:0] down_25_write_in;
  wire down_25_write_write_en;
  wire down_25_write_clk;
  wire [31:0] down_25_write_out;
  wire down_25_write_done;
  wire [31:0] right_25_write_in;
  wire right_25_write_write_en;
  wire right_25_write_clk;
  wire [31:0] right_25_write_out;
  wire right_25_write_done;
  wire [31:0] left_25_read_in;
  wire left_25_read_write_en;
  wire left_25_read_clk;
  wire [31:0] left_25_read_out;
  wire left_25_read_done;
  wire [31:0] top_25_read_in;
  wire top_25_read_write_en;
  wire top_25_read_clk;
  wire [31:0] top_25_read_out;
  wire top_25_read_done;
  wire [31:0] pe_25_top;
  wire [31:0] pe_25_left;
  wire pe_25_go;
  wire pe_25_clk;
  wire [31:0] pe_25_down;
  wire [31:0] pe_25_right;
  wire [31:0] pe_25_out;
  wire pe_25_done;
  wire [31:0] down_24_write_in;
  wire down_24_write_write_en;
  wire down_24_write_clk;
  wire [31:0] down_24_write_out;
  wire down_24_write_done;
  wire [31:0] right_24_write_in;
  wire right_24_write_write_en;
  wire right_24_write_clk;
  wire [31:0] right_24_write_out;
  wire right_24_write_done;
  wire [31:0] left_24_read_in;
  wire left_24_read_write_en;
  wire left_24_read_clk;
  wire [31:0] left_24_read_out;
  wire left_24_read_done;
  wire [31:0] top_24_read_in;
  wire top_24_read_write_en;
  wire top_24_read_clk;
  wire [31:0] top_24_read_out;
  wire top_24_read_done;
  wire [31:0] pe_24_top;
  wire [31:0] pe_24_left;
  wire pe_24_go;
  wire pe_24_clk;
  wire [31:0] pe_24_down;
  wire [31:0] pe_24_right;
  wire [31:0] pe_24_out;
  wire pe_24_done;
  wire [31:0] down_23_write_in;
  wire down_23_write_write_en;
  wire down_23_write_clk;
  wire [31:0] down_23_write_out;
  wire down_23_write_done;
  wire [31:0] right_23_write_in;
  wire right_23_write_write_en;
  wire right_23_write_clk;
  wire [31:0] right_23_write_out;
  wire right_23_write_done;
  wire [31:0] left_23_read_in;
  wire left_23_read_write_en;
  wire left_23_read_clk;
  wire [31:0] left_23_read_out;
  wire left_23_read_done;
  wire [31:0] top_23_read_in;
  wire top_23_read_write_en;
  wire top_23_read_clk;
  wire [31:0] top_23_read_out;
  wire top_23_read_done;
  wire [31:0] pe_23_top;
  wire [31:0] pe_23_left;
  wire pe_23_go;
  wire pe_23_clk;
  wire [31:0] pe_23_down;
  wire [31:0] pe_23_right;
  wire [31:0] pe_23_out;
  wire pe_23_done;
  wire [31:0] down_22_write_in;
  wire down_22_write_write_en;
  wire down_22_write_clk;
  wire [31:0] down_22_write_out;
  wire down_22_write_done;
  wire [31:0] right_22_write_in;
  wire right_22_write_write_en;
  wire right_22_write_clk;
  wire [31:0] right_22_write_out;
  wire right_22_write_done;
  wire [31:0] left_22_read_in;
  wire left_22_read_write_en;
  wire left_22_read_clk;
  wire [31:0] left_22_read_out;
  wire left_22_read_done;
  wire [31:0] top_22_read_in;
  wire top_22_read_write_en;
  wire top_22_read_clk;
  wire [31:0] top_22_read_out;
  wire top_22_read_done;
  wire [31:0] pe_22_top;
  wire [31:0] pe_22_left;
  wire pe_22_go;
  wire pe_22_clk;
  wire [31:0] pe_22_down;
  wire [31:0] pe_22_right;
  wire [31:0] pe_22_out;
  wire pe_22_done;
  wire [31:0] down_21_write_in;
  wire down_21_write_write_en;
  wire down_21_write_clk;
  wire [31:0] down_21_write_out;
  wire down_21_write_done;
  wire [31:0] right_21_write_in;
  wire right_21_write_write_en;
  wire right_21_write_clk;
  wire [31:0] right_21_write_out;
  wire right_21_write_done;
  wire [31:0] left_21_read_in;
  wire left_21_read_write_en;
  wire left_21_read_clk;
  wire [31:0] left_21_read_out;
  wire left_21_read_done;
  wire [31:0] top_21_read_in;
  wire top_21_read_write_en;
  wire top_21_read_clk;
  wire [31:0] top_21_read_out;
  wire top_21_read_done;
  wire [31:0] pe_21_top;
  wire [31:0] pe_21_left;
  wire pe_21_go;
  wire pe_21_clk;
  wire [31:0] pe_21_down;
  wire [31:0] pe_21_right;
  wire [31:0] pe_21_out;
  wire pe_21_done;
  wire [31:0] down_20_write_in;
  wire down_20_write_write_en;
  wire down_20_write_clk;
  wire [31:0] down_20_write_out;
  wire down_20_write_done;
  wire [31:0] right_20_write_in;
  wire right_20_write_write_en;
  wire right_20_write_clk;
  wire [31:0] right_20_write_out;
  wire right_20_write_done;
  wire [31:0] left_20_read_in;
  wire left_20_read_write_en;
  wire left_20_read_clk;
  wire [31:0] left_20_read_out;
  wire left_20_read_done;
  wire [31:0] top_20_read_in;
  wire top_20_read_write_en;
  wire top_20_read_clk;
  wire [31:0] top_20_read_out;
  wire top_20_read_done;
  wire [31:0] pe_20_top;
  wire [31:0] pe_20_left;
  wire pe_20_go;
  wire pe_20_clk;
  wire [31:0] pe_20_down;
  wire [31:0] pe_20_right;
  wire [31:0] pe_20_out;
  wire pe_20_done;
  wire [31:0] down_17_write_in;
  wire down_17_write_write_en;
  wire down_17_write_clk;
  wire [31:0] down_17_write_out;
  wire down_17_write_done;
  wire [31:0] left_17_read_in;
  wire left_17_read_write_en;
  wire left_17_read_clk;
  wire [31:0] left_17_read_out;
  wire left_17_read_done;
  wire [31:0] top_17_read_in;
  wire top_17_read_write_en;
  wire top_17_read_clk;
  wire [31:0] top_17_read_out;
  wire top_17_read_done;
  wire [31:0] pe_17_top;
  wire [31:0] pe_17_left;
  wire pe_17_go;
  wire pe_17_clk;
  wire [31:0] pe_17_down;
  wire [31:0] pe_17_right;
  wire [31:0] pe_17_out;
  wire pe_17_done;
  wire [31:0] down_16_write_in;
  wire down_16_write_write_en;
  wire down_16_write_clk;
  wire [31:0] down_16_write_out;
  wire down_16_write_done;
  wire [31:0] right_16_write_in;
  wire right_16_write_write_en;
  wire right_16_write_clk;
  wire [31:0] right_16_write_out;
  wire right_16_write_done;
  wire [31:0] left_16_read_in;
  wire left_16_read_write_en;
  wire left_16_read_clk;
  wire [31:0] left_16_read_out;
  wire left_16_read_done;
  wire [31:0] top_16_read_in;
  wire top_16_read_write_en;
  wire top_16_read_clk;
  wire [31:0] top_16_read_out;
  wire top_16_read_done;
  wire [31:0] pe_16_top;
  wire [31:0] pe_16_left;
  wire pe_16_go;
  wire pe_16_clk;
  wire [31:0] pe_16_down;
  wire [31:0] pe_16_right;
  wire [31:0] pe_16_out;
  wire pe_16_done;
  wire [31:0] down_15_write_in;
  wire down_15_write_write_en;
  wire down_15_write_clk;
  wire [31:0] down_15_write_out;
  wire down_15_write_done;
  wire [31:0] right_15_write_in;
  wire right_15_write_write_en;
  wire right_15_write_clk;
  wire [31:0] right_15_write_out;
  wire right_15_write_done;
  wire [31:0] left_15_read_in;
  wire left_15_read_write_en;
  wire left_15_read_clk;
  wire [31:0] left_15_read_out;
  wire left_15_read_done;
  wire [31:0] top_15_read_in;
  wire top_15_read_write_en;
  wire top_15_read_clk;
  wire [31:0] top_15_read_out;
  wire top_15_read_done;
  wire [31:0] pe_15_top;
  wire [31:0] pe_15_left;
  wire pe_15_go;
  wire pe_15_clk;
  wire [31:0] pe_15_down;
  wire [31:0] pe_15_right;
  wire [31:0] pe_15_out;
  wire pe_15_done;
  wire [31:0] down_14_write_in;
  wire down_14_write_write_en;
  wire down_14_write_clk;
  wire [31:0] down_14_write_out;
  wire down_14_write_done;
  wire [31:0] right_14_write_in;
  wire right_14_write_write_en;
  wire right_14_write_clk;
  wire [31:0] right_14_write_out;
  wire right_14_write_done;
  wire [31:0] left_14_read_in;
  wire left_14_read_write_en;
  wire left_14_read_clk;
  wire [31:0] left_14_read_out;
  wire left_14_read_done;
  wire [31:0] top_14_read_in;
  wire top_14_read_write_en;
  wire top_14_read_clk;
  wire [31:0] top_14_read_out;
  wire top_14_read_done;
  wire [31:0] pe_14_top;
  wire [31:0] pe_14_left;
  wire pe_14_go;
  wire pe_14_clk;
  wire [31:0] pe_14_down;
  wire [31:0] pe_14_right;
  wire [31:0] pe_14_out;
  wire pe_14_done;
  wire [31:0] down_13_write_in;
  wire down_13_write_write_en;
  wire down_13_write_clk;
  wire [31:0] down_13_write_out;
  wire down_13_write_done;
  wire [31:0] right_13_write_in;
  wire right_13_write_write_en;
  wire right_13_write_clk;
  wire [31:0] right_13_write_out;
  wire right_13_write_done;
  wire [31:0] left_13_read_in;
  wire left_13_read_write_en;
  wire left_13_read_clk;
  wire [31:0] left_13_read_out;
  wire left_13_read_done;
  wire [31:0] top_13_read_in;
  wire top_13_read_write_en;
  wire top_13_read_clk;
  wire [31:0] top_13_read_out;
  wire top_13_read_done;
  wire [31:0] pe_13_top;
  wire [31:0] pe_13_left;
  wire pe_13_go;
  wire pe_13_clk;
  wire [31:0] pe_13_down;
  wire [31:0] pe_13_right;
  wire [31:0] pe_13_out;
  wire pe_13_done;
  wire [31:0] down_12_write_in;
  wire down_12_write_write_en;
  wire down_12_write_clk;
  wire [31:0] down_12_write_out;
  wire down_12_write_done;
  wire [31:0] right_12_write_in;
  wire right_12_write_write_en;
  wire right_12_write_clk;
  wire [31:0] right_12_write_out;
  wire right_12_write_done;
  wire [31:0] left_12_read_in;
  wire left_12_read_write_en;
  wire left_12_read_clk;
  wire [31:0] left_12_read_out;
  wire left_12_read_done;
  wire [31:0] top_12_read_in;
  wire top_12_read_write_en;
  wire top_12_read_clk;
  wire [31:0] top_12_read_out;
  wire top_12_read_done;
  wire [31:0] pe_12_top;
  wire [31:0] pe_12_left;
  wire pe_12_go;
  wire pe_12_clk;
  wire [31:0] pe_12_down;
  wire [31:0] pe_12_right;
  wire [31:0] pe_12_out;
  wire pe_12_done;
  wire [31:0] down_11_write_in;
  wire down_11_write_write_en;
  wire down_11_write_clk;
  wire [31:0] down_11_write_out;
  wire down_11_write_done;
  wire [31:0] right_11_write_in;
  wire right_11_write_write_en;
  wire right_11_write_clk;
  wire [31:0] right_11_write_out;
  wire right_11_write_done;
  wire [31:0] left_11_read_in;
  wire left_11_read_write_en;
  wire left_11_read_clk;
  wire [31:0] left_11_read_out;
  wire left_11_read_done;
  wire [31:0] top_11_read_in;
  wire top_11_read_write_en;
  wire top_11_read_clk;
  wire [31:0] top_11_read_out;
  wire top_11_read_done;
  wire [31:0] pe_11_top;
  wire [31:0] pe_11_left;
  wire pe_11_go;
  wire pe_11_clk;
  wire [31:0] pe_11_down;
  wire [31:0] pe_11_right;
  wire [31:0] pe_11_out;
  wire pe_11_done;
  wire [31:0] down_10_write_in;
  wire down_10_write_write_en;
  wire down_10_write_clk;
  wire [31:0] down_10_write_out;
  wire down_10_write_done;
  wire [31:0] right_10_write_in;
  wire right_10_write_write_en;
  wire right_10_write_clk;
  wire [31:0] right_10_write_out;
  wire right_10_write_done;
  wire [31:0] left_10_read_in;
  wire left_10_read_write_en;
  wire left_10_read_clk;
  wire [31:0] left_10_read_out;
  wire left_10_read_done;
  wire [31:0] top_10_read_in;
  wire top_10_read_write_en;
  wire top_10_read_clk;
  wire [31:0] top_10_read_out;
  wire top_10_read_done;
  wire [31:0] pe_10_top;
  wire [31:0] pe_10_left;
  wire pe_10_go;
  wire pe_10_clk;
  wire [31:0] pe_10_down;
  wire [31:0] pe_10_right;
  wire [31:0] pe_10_out;
  wire pe_10_done;
  wire [31:0] down_07_write_in;
  wire down_07_write_write_en;
  wire down_07_write_clk;
  wire [31:0] down_07_write_out;
  wire down_07_write_done;
  wire [31:0] left_07_read_in;
  wire left_07_read_write_en;
  wire left_07_read_clk;
  wire [31:0] left_07_read_out;
  wire left_07_read_done;
  wire [31:0] top_07_read_in;
  wire top_07_read_write_en;
  wire top_07_read_clk;
  wire [31:0] top_07_read_out;
  wire top_07_read_done;
  wire [31:0] pe_07_top;
  wire [31:0] pe_07_left;
  wire pe_07_go;
  wire pe_07_clk;
  wire [31:0] pe_07_down;
  wire [31:0] pe_07_right;
  wire [31:0] pe_07_out;
  wire pe_07_done;
  wire [31:0] down_06_write_in;
  wire down_06_write_write_en;
  wire down_06_write_clk;
  wire [31:0] down_06_write_out;
  wire down_06_write_done;
  wire [31:0] right_06_write_in;
  wire right_06_write_write_en;
  wire right_06_write_clk;
  wire [31:0] right_06_write_out;
  wire right_06_write_done;
  wire [31:0] left_06_read_in;
  wire left_06_read_write_en;
  wire left_06_read_clk;
  wire [31:0] left_06_read_out;
  wire left_06_read_done;
  wire [31:0] top_06_read_in;
  wire top_06_read_write_en;
  wire top_06_read_clk;
  wire [31:0] top_06_read_out;
  wire top_06_read_done;
  wire [31:0] pe_06_top;
  wire [31:0] pe_06_left;
  wire pe_06_go;
  wire pe_06_clk;
  wire [31:0] pe_06_down;
  wire [31:0] pe_06_right;
  wire [31:0] pe_06_out;
  wire pe_06_done;
  wire [31:0] down_05_write_in;
  wire down_05_write_write_en;
  wire down_05_write_clk;
  wire [31:0] down_05_write_out;
  wire down_05_write_done;
  wire [31:0] right_05_write_in;
  wire right_05_write_write_en;
  wire right_05_write_clk;
  wire [31:0] right_05_write_out;
  wire right_05_write_done;
  wire [31:0] left_05_read_in;
  wire left_05_read_write_en;
  wire left_05_read_clk;
  wire [31:0] left_05_read_out;
  wire left_05_read_done;
  wire [31:0] top_05_read_in;
  wire top_05_read_write_en;
  wire top_05_read_clk;
  wire [31:0] top_05_read_out;
  wire top_05_read_done;
  wire [31:0] pe_05_top;
  wire [31:0] pe_05_left;
  wire pe_05_go;
  wire pe_05_clk;
  wire [31:0] pe_05_down;
  wire [31:0] pe_05_right;
  wire [31:0] pe_05_out;
  wire pe_05_done;
  wire [31:0] down_04_write_in;
  wire down_04_write_write_en;
  wire down_04_write_clk;
  wire [31:0] down_04_write_out;
  wire down_04_write_done;
  wire [31:0] right_04_write_in;
  wire right_04_write_write_en;
  wire right_04_write_clk;
  wire [31:0] right_04_write_out;
  wire right_04_write_done;
  wire [31:0] left_04_read_in;
  wire left_04_read_write_en;
  wire left_04_read_clk;
  wire [31:0] left_04_read_out;
  wire left_04_read_done;
  wire [31:0] top_04_read_in;
  wire top_04_read_write_en;
  wire top_04_read_clk;
  wire [31:0] top_04_read_out;
  wire top_04_read_done;
  wire [31:0] pe_04_top;
  wire [31:0] pe_04_left;
  wire pe_04_go;
  wire pe_04_clk;
  wire [31:0] pe_04_down;
  wire [31:0] pe_04_right;
  wire [31:0] pe_04_out;
  wire pe_04_done;
  wire [31:0] down_03_write_in;
  wire down_03_write_write_en;
  wire down_03_write_clk;
  wire [31:0] down_03_write_out;
  wire down_03_write_done;
  wire [31:0] right_03_write_in;
  wire right_03_write_write_en;
  wire right_03_write_clk;
  wire [31:0] right_03_write_out;
  wire right_03_write_done;
  wire [31:0] left_03_read_in;
  wire left_03_read_write_en;
  wire left_03_read_clk;
  wire [31:0] left_03_read_out;
  wire left_03_read_done;
  wire [31:0] top_03_read_in;
  wire top_03_read_write_en;
  wire top_03_read_clk;
  wire [31:0] top_03_read_out;
  wire top_03_read_done;
  wire [31:0] pe_03_top;
  wire [31:0] pe_03_left;
  wire pe_03_go;
  wire pe_03_clk;
  wire [31:0] pe_03_down;
  wire [31:0] pe_03_right;
  wire [31:0] pe_03_out;
  wire pe_03_done;
  wire [31:0] down_02_write_in;
  wire down_02_write_write_en;
  wire down_02_write_clk;
  wire [31:0] down_02_write_out;
  wire down_02_write_done;
  wire [31:0] right_02_write_in;
  wire right_02_write_write_en;
  wire right_02_write_clk;
  wire [31:0] right_02_write_out;
  wire right_02_write_done;
  wire [31:0] left_02_read_in;
  wire left_02_read_write_en;
  wire left_02_read_clk;
  wire [31:0] left_02_read_out;
  wire left_02_read_done;
  wire [31:0] top_02_read_in;
  wire top_02_read_write_en;
  wire top_02_read_clk;
  wire [31:0] top_02_read_out;
  wire top_02_read_done;
  wire [31:0] pe_02_top;
  wire [31:0] pe_02_left;
  wire pe_02_go;
  wire pe_02_clk;
  wire [31:0] pe_02_down;
  wire [31:0] pe_02_right;
  wire [31:0] pe_02_out;
  wire pe_02_done;
  wire [31:0] down_01_write_in;
  wire down_01_write_write_en;
  wire down_01_write_clk;
  wire [31:0] down_01_write_out;
  wire down_01_write_done;
  wire [31:0] right_01_write_in;
  wire right_01_write_write_en;
  wire right_01_write_clk;
  wire [31:0] right_01_write_out;
  wire right_01_write_done;
  wire [31:0] left_01_read_in;
  wire left_01_read_write_en;
  wire left_01_read_clk;
  wire [31:0] left_01_read_out;
  wire left_01_read_done;
  wire [31:0] top_01_read_in;
  wire top_01_read_write_en;
  wire top_01_read_clk;
  wire [31:0] top_01_read_out;
  wire top_01_read_done;
  wire [31:0] pe_01_top;
  wire [31:0] pe_01_left;
  wire pe_01_go;
  wire pe_01_clk;
  wire [31:0] pe_01_down;
  wire [31:0] pe_01_right;
  wire [31:0] pe_01_out;
  wire pe_01_done;
  wire [31:0] down_00_write_in;
  wire down_00_write_write_en;
  wire down_00_write_clk;
  wire [31:0] down_00_write_out;
  wire down_00_write_done;
  wire [31:0] right_00_write_in;
  wire right_00_write_write_en;
  wire right_00_write_clk;
  wire [31:0] right_00_write_out;
  wire right_00_write_done;
  wire [31:0] left_00_read_in;
  wire left_00_read_write_en;
  wire left_00_read_clk;
  wire [31:0] left_00_read_out;
  wire left_00_read_done;
  wire [31:0] top_00_read_in;
  wire top_00_read_write_en;
  wire top_00_read_clk;
  wire [31:0] top_00_read_out;
  wire top_00_read_done;
  wire [31:0] pe_00_top;
  wire [31:0] pe_00_left;
  wire pe_00_go;
  wire pe_00_clk;
  wire [31:0] pe_00_down;
  wire [31:0] pe_00_right;
  wire [31:0] pe_00_out;
  wire pe_00_done;
  wire [3:0] l7_addr0;
  wire [31:0] l7_write_data;
  wire l7_write_en;
  wire l7_clk;
  wire [31:0] l7_read_data;
  wire l7_done;
  wire [3:0] l7_add_left;
  wire [3:0] l7_add_right;
  wire [3:0] l7_add_out;
  wire [3:0] l7_idx_in;
  wire l7_idx_write_en;
  wire l7_idx_clk;
  wire [3:0] l7_idx_out;
  wire l7_idx_done;
  wire [3:0] l6_addr0;
  wire [31:0] l6_write_data;
  wire l6_write_en;
  wire l6_clk;
  wire [31:0] l6_read_data;
  wire l6_done;
  wire [3:0] l6_add_left;
  wire [3:0] l6_add_right;
  wire [3:0] l6_add_out;
  wire [3:0] l6_idx_in;
  wire l6_idx_write_en;
  wire l6_idx_clk;
  wire [3:0] l6_idx_out;
  wire l6_idx_done;
  wire [3:0] l5_addr0;
  wire [31:0] l5_write_data;
  wire l5_write_en;
  wire l5_clk;
  wire [31:0] l5_read_data;
  wire l5_done;
  wire [3:0] l5_add_left;
  wire [3:0] l5_add_right;
  wire [3:0] l5_add_out;
  wire [3:0] l5_idx_in;
  wire l5_idx_write_en;
  wire l5_idx_clk;
  wire [3:0] l5_idx_out;
  wire l5_idx_done;
  wire [3:0] l4_addr0;
  wire [31:0] l4_write_data;
  wire l4_write_en;
  wire l4_clk;
  wire [31:0] l4_read_data;
  wire l4_done;
  wire [3:0] l4_add_left;
  wire [3:0] l4_add_right;
  wire [3:0] l4_add_out;
  wire [3:0] l4_idx_in;
  wire l4_idx_write_en;
  wire l4_idx_clk;
  wire [3:0] l4_idx_out;
  wire l4_idx_done;
  wire [3:0] l3_addr0;
  wire [31:0] l3_write_data;
  wire l3_write_en;
  wire l3_clk;
  wire [31:0] l3_read_data;
  wire l3_done;
  wire [3:0] l3_add_left;
  wire [3:0] l3_add_right;
  wire [3:0] l3_add_out;
  wire [3:0] l3_idx_in;
  wire l3_idx_write_en;
  wire l3_idx_clk;
  wire [3:0] l3_idx_out;
  wire l3_idx_done;
  wire [3:0] l2_addr0;
  wire [31:0] l2_write_data;
  wire l2_write_en;
  wire l2_clk;
  wire [31:0] l2_read_data;
  wire l2_done;
  wire [3:0] l2_add_left;
  wire [3:0] l2_add_right;
  wire [3:0] l2_add_out;
  wire [3:0] l2_idx_in;
  wire l2_idx_write_en;
  wire l2_idx_clk;
  wire [3:0] l2_idx_out;
  wire l2_idx_done;
  wire [3:0] l1_addr0;
  wire [31:0] l1_write_data;
  wire l1_write_en;
  wire l1_clk;
  wire [31:0] l1_read_data;
  wire l1_done;
  wire [3:0] l1_add_left;
  wire [3:0] l1_add_right;
  wire [3:0] l1_add_out;
  wire [3:0] l1_idx_in;
  wire l1_idx_write_en;
  wire l1_idx_clk;
  wire [3:0] l1_idx_out;
  wire l1_idx_done;
  wire [3:0] l0_addr0;
  wire [31:0] l0_write_data;
  wire l0_write_en;
  wire l0_clk;
  wire [31:0] l0_read_data;
  wire l0_done;
  wire [3:0] l0_add_left;
  wire [3:0] l0_add_right;
  wire [3:0] l0_add_out;
  wire [3:0] l0_idx_in;
  wire l0_idx_write_en;
  wire l0_idx_clk;
  wire [3:0] l0_idx_out;
  wire l0_idx_done;
  wire [3:0] t7_addr0;
  wire [31:0] t7_write_data;
  wire t7_write_en;
  wire t7_clk;
  wire [31:0] t7_read_data;
  wire t7_done;
  wire [3:0] t7_add_left;
  wire [3:0] t7_add_right;
  wire [3:0] t7_add_out;
  wire [3:0] t7_idx_in;
  wire t7_idx_write_en;
  wire t7_idx_clk;
  wire [3:0] t7_idx_out;
  wire t7_idx_done;
  wire [3:0] t6_addr0;
  wire [31:0] t6_write_data;
  wire t6_write_en;
  wire t6_clk;
  wire [31:0] t6_read_data;
  wire t6_done;
  wire [3:0] t6_add_left;
  wire [3:0] t6_add_right;
  wire [3:0] t6_add_out;
  wire [3:0] t6_idx_in;
  wire t6_idx_write_en;
  wire t6_idx_clk;
  wire [3:0] t6_idx_out;
  wire t6_idx_done;
  wire [3:0] t5_addr0;
  wire [31:0] t5_write_data;
  wire t5_write_en;
  wire t5_clk;
  wire [31:0] t5_read_data;
  wire t5_done;
  wire [3:0] t5_add_left;
  wire [3:0] t5_add_right;
  wire [3:0] t5_add_out;
  wire [3:0] t5_idx_in;
  wire t5_idx_write_en;
  wire t5_idx_clk;
  wire [3:0] t5_idx_out;
  wire t5_idx_done;
  wire [3:0] t4_addr0;
  wire [31:0] t4_write_data;
  wire t4_write_en;
  wire t4_clk;
  wire [31:0] t4_read_data;
  wire t4_done;
  wire [3:0] t4_add_left;
  wire [3:0] t4_add_right;
  wire [3:0] t4_add_out;
  wire [3:0] t4_idx_in;
  wire t4_idx_write_en;
  wire t4_idx_clk;
  wire [3:0] t4_idx_out;
  wire t4_idx_done;
  wire [3:0] t3_addr0;
  wire [31:0] t3_write_data;
  wire t3_write_en;
  wire t3_clk;
  wire [31:0] t3_read_data;
  wire t3_done;
  wire [3:0] t3_add_left;
  wire [3:0] t3_add_right;
  wire [3:0] t3_add_out;
  wire [3:0] t3_idx_in;
  wire t3_idx_write_en;
  wire t3_idx_clk;
  wire [3:0] t3_idx_out;
  wire t3_idx_done;
  wire [3:0] t2_addr0;
  wire [31:0] t2_write_data;
  wire t2_write_en;
  wire t2_clk;
  wire [31:0] t2_read_data;
  wire t2_done;
  wire [3:0] t2_add_left;
  wire [3:0] t2_add_right;
  wire [3:0] t2_add_out;
  wire [3:0] t2_idx_in;
  wire t2_idx_write_en;
  wire t2_idx_clk;
  wire [3:0] t2_idx_out;
  wire t2_idx_done;
  wire [3:0] t1_addr0;
  wire [31:0] t1_write_data;
  wire t1_write_en;
  wire t1_clk;
  wire [31:0] t1_read_data;
  wire t1_done;
  wire [3:0] t1_add_left;
  wire [3:0] t1_add_right;
  wire [3:0] t1_add_out;
  wire [3:0] t1_idx_in;
  wire t1_idx_write_en;
  wire t1_idx_clk;
  wire [3:0] t1_idx_out;
  wire t1_idx_done;
  wire [3:0] t0_addr0;
  wire [31:0] t0_write_data;
  wire t0_write_en;
  wire t0_clk;
  wire [31:0] t0_read_data;
  wire t0_done;
  wire [3:0] t0_add_left;
  wire [3:0] t0_add_right;
  wire [3:0] t0_add_out;
  wire [3:0] t0_idx_in;
  wire t0_idx_write_en;
  wire t0_idx_clk;
  wire [3:0] t0_idx_out;
  wire t0_idx_done;
  wire par_reset0_in;
  wire par_reset0_write_en;
  wire par_reset0_clk;
  wire par_reset0_out;
  wire par_reset0_done;
  wire par_done_reg0_in;
  wire par_done_reg0_write_en;
  wire par_done_reg0_clk;
  wire par_done_reg0_out;
  wire par_done_reg0_done;
  wire par_done_reg1_in;
  wire par_done_reg1_write_en;
  wire par_done_reg1_clk;
  wire par_done_reg1_out;
  wire par_done_reg1_done;
  wire par_done_reg2_in;
  wire par_done_reg2_write_en;
  wire par_done_reg2_clk;
  wire par_done_reg2_out;
  wire par_done_reg2_done;
  wire par_done_reg3_in;
  wire par_done_reg3_write_en;
  wire par_done_reg3_clk;
  wire par_done_reg3_out;
  wire par_done_reg3_done;
  wire par_done_reg4_in;
  wire par_done_reg4_write_en;
  wire par_done_reg4_clk;
  wire par_done_reg4_out;
  wire par_done_reg4_done;
  wire par_done_reg5_in;
  wire par_done_reg5_write_en;
  wire par_done_reg5_clk;
  wire par_done_reg5_out;
  wire par_done_reg5_done;
  wire par_done_reg6_in;
  wire par_done_reg6_write_en;
  wire par_done_reg6_clk;
  wire par_done_reg6_out;
  wire par_done_reg6_done;
  wire par_done_reg7_in;
  wire par_done_reg7_write_en;
  wire par_done_reg7_clk;
  wire par_done_reg7_out;
  wire par_done_reg7_done;
  wire par_done_reg8_in;
  wire par_done_reg8_write_en;
  wire par_done_reg8_clk;
  wire par_done_reg8_out;
  wire par_done_reg8_done;
  wire par_done_reg9_in;
  wire par_done_reg9_write_en;
  wire par_done_reg9_clk;
  wire par_done_reg9_out;
  wire par_done_reg9_done;
  wire par_done_reg10_in;
  wire par_done_reg10_write_en;
  wire par_done_reg10_clk;
  wire par_done_reg10_out;
  wire par_done_reg10_done;
  wire par_done_reg11_in;
  wire par_done_reg11_write_en;
  wire par_done_reg11_clk;
  wire par_done_reg11_out;
  wire par_done_reg11_done;
  wire par_done_reg12_in;
  wire par_done_reg12_write_en;
  wire par_done_reg12_clk;
  wire par_done_reg12_out;
  wire par_done_reg12_done;
  wire par_done_reg13_in;
  wire par_done_reg13_write_en;
  wire par_done_reg13_clk;
  wire par_done_reg13_out;
  wire par_done_reg13_done;
  wire par_done_reg14_in;
  wire par_done_reg14_write_en;
  wire par_done_reg14_clk;
  wire par_done_reg14_out;
  wire par_done_reg14_done;
  wire par_done_reg15_in;
  wire par_done_reg15_write_en;
  wire par_done_reg15_clk;
  wire par_done_reg15_out;
  wire par_done_reg15_done;
  wire par_reset1_in;
  wire par_reset1_write_en;
  wire par_reset1_clk;
  wire par_reset1_out;
  wire par_reset1_done;
  wire par_done_reg16_in;
  wire par_done_reg16_write_en;
  wire par_done_reg16_clk;
  wire par_done_reg16_out;
  wire par_done_reg16_done;
  wire par_done_reg17_in;
  wire par_done_reg17_write_en;
  wire par_done_reg17_clk;
  wire par_done_reg17_out;
  wire par_done_reg17_done;
  wire par_reset2_in;
  wire par_reset2_write_en;
  wire par_reset2_clk;
  wire par_reset2_out;
  wire par_reset2_done;
  wire par_done_reg18_in;
  wire par_done_reg18_write_en;
  wire par_done_reg18_clk;
  wire par_done_reg18_out;
  wire par_done_reg18_done;
  wire par_done_reg19_in;
  wire par_done_reg19_write_en;
  wire par_done_reg19_clk;
  wire par_done_reg19_out;
  wire par_done_reg19_done;
  wire par_reset3_in;
  wire par_reset3_write_en;
  wire par_reset3_clk;
  wire par_reset3_out;
  wire par_reset3_done;
  wire par_done_reg20_in;
  wire par_done_reg20_write_en;
  wire par_done_reg20_clk;
  wire par_done_reg20_out;
  wire par_done_reg20_done;
  wire par_done_reg21_in;
  wire par_done_reg21_write_en;
  wire par_done_reg21_clk;
  wire par_done_reg21_out;
  wire par_done_reg21_done;
  wire par_done_reg22_in;
  wire par_done_reg22_write_en;
  wire par_done_reg22_clk;
  wire par_done_reg22_out;
  wire par_done_reg22_done;
  wire par_done_reg23_in;
  wire par_done_reg23_write_en;
  wire par_done_reg23_clk;
  wire par_done_reg23_out;
  wire par_done_reg23_done;
  wire par_done_reg24_in;
  wire par_done_reg24_write_en;
  wire par_done_reg24_clk;
  wire par_done_reg24_out;
  wire par_done_reg24_done;
  wire par_reset4_in;
  wire par_reset4_write_en;
  wire par_reset4_clk;
  wire par_reset4_out;
  wire par_reset4_done;
  wire par_done_reg25_in;
  wire par_done_reg25_write_en;
  wire par_done_reg25_clk;
  wire par_done_reg25_out;
  wire par_done_reg25_done;
  wire par_done_reg26_in;
  wire par_done_reg26_write_en;
  wire par_done_reg26_clk;
  wire par_done_reg26_out;
  wire par_done_reg26_done;
  wire par_done_reg27_in;
  wire par_done_reg27_write_en;
  wire par_done_reg27_clk;
  wire par_done_reg27_out;
  wire par_done_reg27_done;
  wire par_done_reg28_in;
  wire par_done_reg28_write_en;
  wire par_done_reg28_clk;
  wire par_done_reg28_out;
  wire par_done_reg28_done;
  wire par_done_reg29_in;
  wire par_done_reg29_write_en;
  wire par_done_reg29_clk;
  wire par_done_reg29_out;
  wire par_done_reg29_done;
  wire par_done_reg30_in;
  wire par_done_reg30_write_en;
  wire par_done_reg30_clk;
  wire par_done_reg30_out;
  wire par_done_reg30_done;
  wire par_reset5_in;
  wire par_reset5_write_en;
  wire par_reset5_clk;
  wire par_reset5_out;
  wire par_reset5_done;
  wire par_done_reg31_in;
  wire par_done_reg31_write_en;
  wire par_done_reg31_clk;
  wire par_done_reg31_out;
  wire par_done_reg31_done;
  wire par_done_reg32_in;
  wire par_done_reg32_write_en;
  wire par_done_reg32_clk;
  wire par_done_reg32_out;
  wire par_done_reg32_done;
  wire par_done_reg33_in;
  wire par_done_reg33_write_en;
  wire par_done_reg33_clk;
  wire par_done_reg33_out;
  wire par_done_reg33_done;
  wire par_done_reg34_in;
  wire par_done_reg34_write_en;
  wire par_done_reg34_clk;
  wire par_done_reg34_out;
  wire par_done_reg34_done;
  wire par_done_reg35_in;
  wire par_done_reg35_write_en;
  wire par_done_reg35_clk;
  wire par_done_reg35_out;
  wire par_done_reg35_done;
  wire par_done_reg36_in;
  wire par_done_reg36_write_en;
  wire par_done_reg36_clk;
  wire par_done_reg36_out;
  wire par_done_reg36_done;
  wire par_done_reg37_in;
  wire par_done_reg37_write_en;
  wire par_done_reg37_clk;
  wire par_done_reg37_out;
  wire par_done_reg37_done;
  wire par_done_reg38_in;
  wire par_done_reg38_write_en;
  wire par_done_reg38_clk;
  wire par_done_reg38_out;
  wire par_done_reg38_done;
  wire par_done_reg39_in;
  wire par_done_reg39_write_en;
  wire par_done_reg39_clk;
  wire par_done_reg39_out;
  wire par_done_reg39_done;
  wire par_reset6_in;
  wire par_reset6_write_en;
  wire par_reset6_clk;
  wire par_reset6_out;
  wire par_reset6_done;
  wire par_done_reg40_in;
  wire par_done_reg40_write_en;
  wire par_done_reg40_clk;
  wire par_done_reg40_out;
  wire par_done_reg40_done;
  wire par_done_reg41_in;
  wire par_done_reg41_write_en;
  wire par_done_reg41_clk;
  wire par_done_reg41_out;
  wire par_done_reg41_done;
  wire par_done_reg42_in;
  wire par_done_reg42_write_en;
  wire par_done_reg42_clk;
  wire par_done_reg42_out;
  wire par_done_reg42_done;
  wire par_done_reg43_in;
  wire par_done_reg43_write_en;
  wire par_done_reg43_clk;
  wire par_done_reg43_out;
  wire par_done_reg43_done;
  wire par_done_reg44_in;
  wire par_done_reg44_write_en;
  wire par_done_reg44_clk;
  wire par_done_reg44_out;
  wire par_done_reg44_done;
  wire par_done_reg45_in;
  wire par_done_reg45_write_en;
  wire par_done_reg45_clk;
  wire par_done_reg45_out;
  wire par_done_reg45_done;
  wire par_done_reg46_in;
  wire par_done_reg46_write_en;
  wire par_done_reg46_clk;
  wire par_done_reg46_out;
  wire par_done_reg46_done;
  wire par_done_reg47_in;
  wire par_done_reg47_write_en;
  wire par_done_reg47_clk;
  wire par_done_reg47_out;
  wire par_done_reg47_done;
  wire par_done_reg48_in;
  wire par_done_reg48_write_en;
  wire par_done_reg48_clk;
  wire par_done_reg48_out;
  wire par_done_reg48_done;
  wire par_done_reg49_in;
  wire par_done_reg49_write_en;
  wire par_done_reg49_clk;
  wire par_done_reg49_out;
  wire par_done_reg49_done;
  wire par_done_reg50_in;
  wire par_done_reg50_write_en;
  wire par_done_reg50_clk;
  wire par_done_reg50_out;
  wire par_done_reg50_done;
  wire par_done_reg51_in;
  wire par_done_reg51_write_en;
  wire par_done_reg51_clk;
  wire par_done_reg51_out;
  wire par_done_reg51_done;
  wire par_reset7_in;
  wire par_reset7_write_en;
  wire par_reset7_clk;
  wire par_reset7_out;
  wire par_reset7_done;
  wire par_done_reg52_in;
  wire par_done_reg52_write_en;
  wire par_done_reg52_clk;
  wire par_done_reg52_out;
  wire par_done_reg52_done;
  wire par_done_reg53_in;
  wire par_done_reg53_write_en;
  wire par_done_reg53_clk;
  wire par_done_reg53_out;
  wire par_done_reg53_done;
  wire par_done_reg54_in;
  wire par_done_reg54_write_en;
  wire par_done_reg54_clk;
  wire par_done_reg54_out;
  wire par_done_reg54_done;
  wire par_done_reg55_in;
  wire par_done_reg55_write_en;
  wire par_done_reg55_clk;
  wire par_done_reg55_out;
  wire par_done_reg55_done;
  wire par_done_reg56_in;
  wire par_done_reg56_write_en;
  wire par_done_reg56_clk;
  wire par_done_reg56_out;
  wire par_done_reg56_done;
  wire par_done_reg57_in;
  wire par_done_reg57_write_en;
  wire par_done_reg57_clk;
  wire par_done_reg57_out;
  wire par_done_reg57_done;
  wire par_done_reg58_in;
  wire par_done_reg58_write_en;
  wire par_done_reg58_clk;
  wire par_done_reg58_out;
  wire par_done_reg58_done;
  wire par_done_reg59_in;
  wire par_done_reg59_write_en;
  wire par_done_reg59_clk;
  wire par_done_reg59_out;
  wire par_done_reg59_done;
  wire par_done_reg60_in;
  wire par_done_reg60_write_en;
  wire par_done_reg60_clk;
  wire par_done_reg60_out;
  wire par_done_reg60_done;
  wire par_done_reg61_in;
  wire par_done_reg61_write_en;
  wire par_done_reg61_clk;
  wire par_done_reg61_out;
  wire par_done_reg61_done;
  wire par_done_reg62_in;
  wire par_done_reg62_write_en;
  wire par_done_reg62_clk;
  wire par_done_reg62_out;
  wire par_done_reg62_done;
  wire par_done_reg63_in;
  wire par_done_reg63_write_en;
  wire par_done_reg63_clk;
  wire par_done_reg63_out;
  wire par_done_reg63_done;
  wire par_done_reg64_in;
  wire par_done_reg64_write_en;
  wire par_done_reg64_clk;
  wire par_done_reg64_out;
  wire par_done_reg64_done;
  wire par_done_reg65_in;
  wire par_done_reg65_write_en;
  wire par_done_reg65_clk;
  wire par_done_reg65_out;
  wire par_done_reg65_done;
  wire par_reset8_in;
  wire par_reset8_write_en;
  wire par_reset8_clk;
  wire par_reset8_out;
  wire par_reset8_done;
  wire par_done_reg66_in;
  wire par_done_reg66_write_en;
  wire par_done_reg66_clk;
  wire par_done_reg66_out;
  wire par_done_reg66_done;
  wire par_done_reg67_in;
  wire par_done_reg67_write_en;
  wire par_done_reg67_clk;
  wire par_done_reg67_out;
  wire par_done_reg67_done;
  wire par_done_reg68_in;
  wire par_done_reg68_write_en;
  wire par_done_reg68_clk;
  wire par_done_reg68_out;
  wire par_done_reg68_done;
  wire par_done_reg69_in;
  wire par_done_reg69_write_en;
  wire par_done_reg69_clk;
  wire par_done_reg69_out;
  wire par_done_reg69_done;
  wire par_done_reg70_in;
  wire par_done_reg70_write_en;
  wire par_done_reg70_clk;
  wire par_done_reg70_out;
  wire par_done_reg70_done;
  wire par_done_reg71_in;
  wire par_done_reg71_write_en;
  wire par_done_reg71_clk;
  wire par_done_reg71_out;
  wire par_done_reg71_done;
  wire par_done_reg72_in;
  wire par_done_reg72_write_en;
  wire par_done_reg72_clk;
  wire par_done_reg72_out;
  wire par_done_reg72_done;
  wire par_done_reg73_in;
  wire par_done_reg73_write_en;
  wire par_done_reg73_clk;
  wire par_done_reg73_out;
  wire par_done_reg73_done;
  wire par_done_reg74_in;
  wire par_done_reg74_write_en;
  wire par_done_reg74_clk;
  wire par_done_reg74_out;
  wire par_done_reg74_done;
  wire par_done_reg75_in;
  wire par_done_reg75_write_en;
  wire par_done_reg75_clk;
  wire par_done_reg75_out;
  wire par_done_reg75_done;
  wire par_done_reg76_in;
  wire par_done_reg76_write_en;
  wire par_done_reg76_clk;
  wire par_done_reg76_out;
  wire par_done_reg76_done;
  wire par_done_reg77_in;
  wire par_done_reg77_write_en;
  wire par_done_reg77_clk;
  wire par_done_reg77_out;
  wire par_done_reg77_done;
  wire par_done_reg78_in;
  wire par_done_reg78_write_en;
  wire par_done_reg78_clk;
  wire par_done_reg78_out;
  wire par_done_reg78_done;
  wire par_done_reg79_in;
  wire par_done_reg79_write_en;
  wire par_done_reg79_clk;
  wire par_done_reg79_out;
  wire par_done_reg79_done;
  wire par_done_reg80_in;
  wire par_done_reg80_write_en;
  wire par_done_reg80_clk;
  wire par_done_reg80_out;
  wire par_done_reg80_done;
  wire par_done_reg81_in;
  wire par_done_reg81_write_en;
  wire par_done_reg81_clk;
  wire par_done_reg81_out;
  wire par_done_reg81_done;
  wire par_done_reg82_in;
  wire par_done_reg82_write_en;
  wire par_done_reg82_clk;
  wire par_done_reg82_out;
  wire par_done_reg82_done;
  wire par_done_reg83_in;
  wire par_done_reg83_write_en;
  wire par_done_reg83_clk;
  wire par_done_reg83_out;
  wire par_done_reg83_done;
  wire par_done_reg84_in;
  wire par_done_reg84_write_en;
  wire par_done_reg84_clk;
  wire par_done_reg84_out;
  wire par_done_reg84_done;
  wire par_done_reg85_in;
  wire par_done_reg85_write_en;
  wire par_done_reg85_clk;
  wire par_done_reg85_out;
  wire par_done_reg85_done;
  wire par_reset9_in;
  wire par_reset9_write_en;
  wire par_reset9_clk;
  wire par_reset9_out;
  wire par_reset9_done;
  wire par_done_reg86_in;
  wire par_done_reg86_write_en;
  wire par_done_reg86_clk;
  wire par_done_reg86_out;
  wire par_done_reg86_done;
  wire par_done_reg87_in;
  wire par_done_reg87_write_en;
  wire par_done_reg87_clk;
  wire par_done_reg87_out;
  wire par_done_reg87_done;
  wire par_done_reg88_in;
  wire par_done_reg88_write_en;
  wire par_done_reg88_clk;
  wire par_done_reg88_out;
  wire par_done_reg88_done;
  wire par_done_reg89_in;
  wire par_done_reg89_write_en;
  wire par_done_reg89_clk;
  wire par_done_reg89_out;
  wire par_done_reg89_done;
  wire par_done_reg90_in;
  wire par_done_reg90_write_en;
  wire par_done_reg90_clk;
  wire par_done_reg90_out;
  wire par_done_reg90_done;
  wire par_done_reg91_in;
  wire par_done_reg91_write_en;
  wire par_done_reg91_clk;
  wire par_done_reg91_out;
  wire par_done_reg91_done;
  wire par_done_reg92_in;
  wire par_done_reg92_write_en;
  wire par_done_reg92_clk;
  wire par_done_reg92_out;
  wire par_done_reg92_done;
  wire par_done_reg93_in;
  wire par_done_reg93_write_en;
  wire par_done_reg93_clk;
  wire par_done_reg93_out;
  wire par_done_reg93_done;
  wire par_done_reg94_in;
  wire par_done_reg94_write_en;
  wire par_done_reg94_clk;
  wire par_done_reg94_out;
  wire par_done_reg94_done;
  wire par_done_reg95_in;
  wire par_done_reg95_write_en;
  wire par_done_reg95_clk;
  wire par_done_reg95_out;
  wire par_done_reg95_done;
  wire par_done_reg96_in;
  wire par_done_reg96_write_en;
  wire par_done_reg96_clk;
  wire par_done_reg96_out;
  wire par_done_reg96_done;
  wire par_done_reg97_in;
  wire par_done_reg97_write_en;
  wire par_done_reg97_clk;
  wire par_done_reg97_out;
  wire par_done_reg97_done;
  wire par_done_reg98_in;
  wire par_done_reg98_write_en;
  wire par_done_reg98_clk;
  wire par_done_reg98_out;
  wire par_done_reg98_done;
  wire par_done_reg99_in;
  wire par_done_reg99_write_en;
  wire par_done_reg99_clk;
  wire par_done_reg99_out;
  wire par_done_reg99_done;
  wire par_done_reg100_in;
  wire par_done_reg100_write_en;
  wire par_done_reg100_clk;
  wire par_done_reg100_out;
  wire par_done_reg100_done;
  wire par_done_reg101_in;
  wire par_done_reg101_write_en;
  wire par_done_reg101_clk;
  wire par_done_reg101_out;
  wire par_done_reg101_done;
  wire par_done_reg102_in;
  wire par_done_reg102_write_en;
  wire par_done_reg102_clk;
  wire par_done_reg102_out;
  wire par_done_reg102_done;
  wire par_done_reg103_in;
  wire par_done_reg103_write_en;
  wire par_done_reg103_clk;
  wire par_done_reg103_out;
  wire par_done_reg103_done;
  wire par_done_reg104_in;
  wire par_done_reg104_write_en;
  wire par_done_reg104_clk;
  wire par_done_reg104_out;
  wire par_done_reg104_done;
  wire par_done_reg105_in;
  wire par_done_reg105_write_en;
  wire par_done_reg105_clk;
  wire par_done_reg105_out;
  wire par_done_reg105_done;
  wire par_reset10_in;
  wire par_reset10_write_en;
  wire par_reset10_clk;
  wire par_reset10_out;
  wire par_reset10_done;
  wire par_done_reg106_in;
  wire par_done_reg106_write_en;
  wire par_done_reg106_clk;
  wire par_done_reg106_out;
  wire par_done_reg106_done;
  wire par_done_reg107_in;
  wire par_done_reg107_write_en;
  wire par_done_reg107_clk;
  wire par_done_reg107_out;
  wire par_done_reg107_done;
  wire par_done_reg108_in;
  wire par_done_reg108_write_en;
  wire par_done_reg108_clk;
  wire par_done_reg108_out;
  wire par_done_reg108_done;
  wire par_done_reg109_in;
  wire par_done_reg109_write_en;
  wire par_done_reg109_clk;
  wire par_done_reg109_out;
  wire par_done_reg109_done;
  wire par_done_reg110_in;
  wire par_done_reg110_write_en;
  wire par_done_reg110_clk;
  wire par_done_reg110_out;
  wire par_done_reg110_done;
  wire par_done_reg111_in;
  wire par_done_reg111_write_en;
  wire par_done_reg111_clk;
  wire par_done_reg111_out;
  wire par_done_reg111_done;
  wire par_done_reg112_in;
  wire par_done_reg112_write_en;
  wire par_done_reg112_clk;
  wire par_done_reg112_out;
  wire par_done_reg112_done;
  wire par_done_reg113_in;
  wire par_done_reg113_write_en;
  wire par_done_reg113_clk;
  wire par_done_reg113_out;
  wire par_done_reg113_done;
  wire par_done_reg114_in;
  wire par_done_reg114_write_en;
  wire par_done_reg114_clk;
  wire par_done_reg114_out;
  wire par_done_reg114_done;
  wire par_done_reg115_in;
  wire par_done_reg115_write_en;
  wire par_done_reg115_clk;
  wire par_done_reg115_out;
  wire par_done_reg115_done;
  wire par_done_reg116_in;
  wire par_done_reg116_write_en;
  wire par_done_reg116_clk;
  wire par_done_reg116_out;
  wire par_done_reg116_done;
  wire par_done_reg117_in;
  wire par_done_reg117_write_en;
  wire par_done_reg117_clk;
  wire par_done_reg117_out;
  wire par_done_reg117_done;
  wire par_done_reg118_in;
  wire par_done_reg118_write_en;
  wire par_done_reg118_clk;
  wire par_done_reg118_out;
  wire par_done_reg118_done;
  wire par_done_reg119_in;
  wire par_done_reg119_write_en;
  wire par_done_reg119_clk;
  wire par_done_reg119_out;
  wire par_done_reg119_done;
  wire par_done_reg120_in;
  wire par_done_reg120_write_en;
  wire par_done_reg120_clk;
  wire par_done_reg120_out;
  wire par_done_reg120_done;
  wire par_done_reg121_in;
  wire par_done_reg121_write_en;
  wire par_done_reg121_clk;
  wire par_done_reg121_out;
  wire par_done_reg121_done;
  wire par_done_reg122_in;
  wire par_done_reg122_write_en;
  wire par_done_reg122_clk;
  wire par_done_reg122_out;
  wire par_done_reg122_done;
  wire par_done_reg123_in;
  wire par_done_reg123_write_en;
  wire par_done_reg123_clk;
  wire par_done_reg123_out;
  wire par_done_reg123_done;
  wire par_done_reg124_in;
  wire par_done_reg124_write_en;
  wire par_done_reg124_clk;
  wire par_done_reg124_out;
  wire par_done_reg124_done;
  wire par_done_reg125_in;
  wire par_done_reg125_write_en;
  wire par_done_reg125_clk;
  wire par_done_reg125_out;
  wire par_done_reg125_done;
  wire par_done_reg126_in;
  wire par_done_reg126_write_en;
  wire par_done_reg126_clk;
  wire par_done_reg126_out;
  wire par_done_reg126_done;
  wire par_done_reg127_in;
  wire par_done_reg127_write_en;
  wire par_done_reg127_clk;
  wire par_done_reg127_out;
  wire par_done_reg127_done;
  wire par_done_reg128_in;
  wire par_done_reg128_write_en;
  wire par_done_reg128_clk;
  wire par_done_reg128_out;
  wire par_done_reg128_done;
  wire par_done_reg129_in;
  wire par_done_reg129_write_en;
  wire par_done_reg129_clk;
  wire par_done_reg129_out;
  wire par_done_reg129_done;
  wire par_done_reg130_in;
  wire par_done_reg130_write_en;
  wire par_done_reg130_clk;
  wire par_done_reg130_out;
  wire par_done_reg130_done;
  wire par_done_reg131_in;
  wire par_done_reg131_write_en;
  wire par_done_reg131_clk;
  wire par_done_reg131_out;
  wire par_done_reg131_done;
  wire par_done_reg132_in;
  wire par_done_reg132_write_en;
  wire par_done_reg132_clk;
  wire par_done_reg132_out;
  wire par_done_reg132_done;
  wire par_done_reg133_in;
  wire par_done_reg133_write_en;
  wire par_done_reg133_clk;
  wire par_done_reg133_out;
  wire par_done_reg133_done;
  wire par_done_reg134_in;
  wire par_done_reg134_write_en;
  wire par_done_reg134_clk;
  wire par_done_reg134_out;
  wire par_done_reg134_done;
  wire par_done_reg135_in;
  wire par_done_reg135_write_en;
  wire par_done_reg135_clk;
  wire par_done_reg135_out;
  wire par_done_reg135_done;
  wire par_reset11_in;
  wire par_reset11_write_en;
  wire par_reset11_clk;
  wire par_reset11_out;
  wire par_reset11_done;
  wire par_done_reg136_in;
  wire par_done_reg136_write_en;
  wire par_done_reg136_clk;
  wire par_done_reg136_out;
  wire par_done_reg136_done;
  wire par_done_reg137_in;
  wire par_done_reg137_write_en;
  wire par_done_reg137_clk;
  wire par_done_reg137_out;
  wire par_done_reg137_done;
  wire par_done_reg138_in;
  wire par_done_reg138_write_en;
  wire par_done_reg138_clk;
  wire par_done_reg138_out;
  wire par_done_reg138_done;
  wire par_done_reg139_in;
  wire par_done_reg139_write_en;
  wire par_done_reg139_clk;
  wire par_done_reg139_out;
  wire par_done_reg139_done;
  wire par_done_reg140_in;
  wire par_done_reg140_write_en;
  wire par_done_reg140_clk;
  wire par_done_reg140_out;
  wire par_done_reg140_done;
  wire par_done_reg141_in;
  wire par_done_reg141_write_en;
  wire par_done_reg141_clk;
  wire par_done_reg141_out;
  wire par_done_reg141_done;
  wire par_done_reg142_in;
  wire par_done_reg142_write_en;
  wire par_done_reg142_clk;
  wire par_done_reg142_out;
  wire par_done_reg142_done;
  wire par_done_reg143_in;
  wire par_done_reg143_write_en;
  wire par_done_reg143_clk;
  wire par_done_reg143_out;
  wire par_done_reg143_done;
  wire par_done_reg144_in;
  wire par_done_reg144_write_en;
  wire par_done_reg144_clk;
  wire par_done_reg144_out;
  wire par_done_reg144_done;
  wire par_done_reg145_in;
  wire par_done_reg145_write_en;
  wire par_done_reg145_clk;
  wire par_done_reg145_out;
  wire par_done_reg145_done;
  wire par_done_reg146_in;
  wire par_done_reg146_write_en;
  wire par_done_reg146_clk;
  wire par_done_reg146_out;
  wire par_done_reg146_done;
  wire par_done_reg147_in;
  wire par_done_reg147_write_en;
  wire par_done_reg147_clk;
  wire par_done_reg147_out;
  wire par_done_reg147_done;
  wire par_done_reg148_in;
  wire par_done_reg148_write_en;
  wire par_done_reg148_clk;
  wire par_done_reg148_out;
  wire par_done_reg148_done;
  wire par_done_reg149_in;
  wire par_done_reg149_write_en;
  wire par_done_reg149_clk;
  wire par_done_reg149_out;
  wire par_done_reg149_done;
  wire par_done_reg150_in;
  wire par_done_reg150_write_en;
  wire par_done_reg150_clk;
  wire par_done_reg150_out;
  wire par_done_reg150_done;
  wire par_done_reg151_in;
  wire par_done_reg151_write_en;
  wire par_done_reg151_clk;
  wire par_done_reg151_out;
  wire par_done_reg151_done;
  wire par_done_reg152_in;
  wire par_done_reg152_write_en;
  wire par_done_reg152_clk;
  wire par_done_reg152_out;
  wire par_done_reg152_done;
  wire par_done_reg153_in;
  wire par_done_reg153_write_en;
  wire par_done_reg153_clk;
  wire par_done_reg153_out;
  wire par_done_reg153_done;
  wire par_done_reg154_in;
  wire par_done_reg154_write_en;
  wire par_done_reg154_clk;
  wire par_done_reg154_out;
  wire par_done_reg154_done;
  wire par_done_reg155_in;
  wire par_done_reg155_write_en;
  wire par_done_reg155_clk;
  wire par_done_reg155_out;
  wire par_done_reg155_done;
  wire par_done_reg156_in;
  wire par_done_reg156_write_en;
  wire par_done_reg156_clk;
  wire par_done_reg156_out;
  wire par_done_reg156_done;
  wire par_done_reg157_in;
  wire par_done_reg157_write_en;
  wire par_done_reg157_clk;
  wire par_done_reg157_out;
  wire par_done_reg157_done;
  wire par_done_reg158_in;
  wire par_done_reg158_write_en;
  wire par_done_reg158_clk;
  wire par_done_reg158_out;
  wire par_done_reg158_done;
  wire par_done_reg159_in;
  wire par_done_reg159_write_en;
  wire par_done_reg159_clk;
  wire par_done_reg159_out;
  wire par_done_reg159_done;
  wire par_done_reg160_in;
  wire par_done_reg160_write_en;
  wire par_done_reg160_clk;
  wire par_done_reg160_out;
  wire par_done_reg160_done;
  wire par_done_reg161_in;
  wire par_done_reg161_write_en;
  wire par_done_reg161_clk;
  wire par_done_reg161_out;
  wire par_done_reg161_done;
  wire par_done_reg162_in;
  wire par_done_reg162_write_en;
  wire par_done_reg162_clk;
  wire par_done_reg162_out;
  wire par_done_reg162_done;
  wire par_reset12_in;
  wire par_reset12_write_en;
  wire par_reset12_clk;
  wire par_reset12_out;
  wire par_reset12_done;
  wire par_done_reg163_in;
  wire par_done_reg163_write_en;
  wire par_done_reg163_clk;
  wire par_done_reg163_out;
  wire par_done_reg163_done;
  wire par_done_reg164_in;
  wire par_done_reg164_write_en;
  wire par_done_reg164_clk;
  wire par_done_reg164_out;
  wire par_done_reg164_done;
  wire par_done_reg165_in;
  wire par_done_reg165_write_en;
  wire par_done_reg165_clk;
  wire par_done_reg165_out;
  wire par_done_reg165_done;
  wire par_done_reg166_in;
  wire par_done_reg166_write_en;
  wire par_done_reg166_clk;
  wire par_done_reg166_out;
  wire par_done_reg166_done;
  wire par_done_reg167_in;
  wire par_done_reg167_write_en;
  wire par_done_reg167_clk;
  wire par_done_reg167_out;
  wire par_done_reg167_done;
  wire par_done_reg168_in;
  wire par_done_reg168_write_en;
  wire par_done_reg168_clk;
  wire par_done_reg168_out;
  wire par_done_reg168_done;
  wire par_done_reg169_in;
  wire par_done_reg169_write_en;
  wire par_done_reg169_clk;
  wire par_done_reg169_out;
  wire par_done_reg169_done;
  wire par_done_reg170_in;
  wire par_done_reg170_write_en;
  wire par_done_reg170_clk;
  wire par_done_reg170_out;
  wire par_done_reg170_done;
  wire par_done_reg171_in;
  wire par_done_reg171_write_en;
  wire par_done_reg171_clk;
  wire par_done_reg171_out;
  wire par_done_reg171_done;
  wire par_done_reg172_in;
  wire par_done_reg172_write_en;
  wire par_done_reg172_clk;
  wire par_done_reg172_out;
  wire par_done_reg172_done;
  wire par_done_reg173_in;
  wire par_done_reg173_write_en;
  wire par_done_reg173_clk;
  wire par_done_reg173_out;
  wire par_done_reg173_done;
  wire par_done_reg174_in;
  wire par_done_reg174_write_en;
  wire par_done_reg174_clk;
  wire par_done_reg174_out;
  wire par_done_reg174_done;
  wire par_done_reg175_in;
  wire par_done_reg175_write_en;
  wire par_done_reg175_clk;
  wire par_done_reg175_out;
  wire par_done_reg175_done;
  wire par_done_reg176_in;
  wire par_done_reg176_write_en;
  wire par_done_reg176_clk;
  wire par_done_reg176_out;
  wire par_done_reg176_done;
  wire par_done_reg177_in;
  wire par_done_reg177_write_en;
  wire par_done_reg177_clk;
  wire par_done_reg177_out;
  wire par_done_reg177_done;
  wire par_done_reg178_in;
  wire par_done_reg178_write_en;
  wire par_done_reg178_clk;
  wire par_done_reg178_out;
  wire par_done_reg178_done;
  wire par_done_reg179_in;
  wire par_done_reg179_write_en;
  wire par_done_reg179_clk;
  wire par_done_reg179_out;
  wire par_done_reg179_done;
  wire par_done_reg180_in;
  wire par_done_reg180_write_en;
  wire par_done_reg180_clk;
  wire par_done_reg180_out;
  wire par_done_reg180_done;
  wire par_done_reg181_in;
  wire par_done_reg181_write_en;
  wire par_done_reg181_clk;
  wire par_done_reg181_out;
  wire par_done_reg181_done;
  wire par_done_reg182_in;
  wire par_done_reg182_write_en;
  wire par_done_reg182_clk;
  wire par_done_reg182_out;
  wire par_done_reg182_done;
  wire par_done_reg183_in;
  wire par_done_reg183_write_en;
  wire par_done_reg183_clk;
  wire par_done_reg183_out;
  wire par_done_reg183_done;
  wire par_done_reg184_in;
  wire par_done_reg184_write_en;
  wire par_done_reg184_clk;
  wire par_done_reg184_out;
  wire par_done_reg184_done;
  wire par_done_reg185_in;
  wire par_done_reg185_write_en;
  wire par_done_reg185_clk;
  wire par_done_reg185_out;
  wire par_done_reg185_done;
  wire par_done_reg186_in;
  wire par_done_reg186_write_en;
  wire par_done_reg186_clk;
  wire par_done_reg186_out;
  wire par_done_reg186_done;
  wire par_done_reg187_in;
  wire par_done_reg187_write_en;
  wire par_done_reg187_clk;
  wire par_done_reg187_out;
  wire par_done_reg187_done;
  wire par_done_reg188_in;
  wire par_done_reg188_write_en;
  wire par_done_reg188_clk;
  wire par_done_reg188_out;
  wire par_done_reg188_done;
  wire par_done_reg189_in;
  wire par_done_reg189_write_en;
  wire par_done_reg189_clk;
  wire par_done_reg189_out;
  wire par_done_reg189_done;
  wire par_done_reg190_in;
  wire par_done_reg190_write_en;
  wire par_done_reg190_clk;
  wire par_done_reg190_out;
  wire par_done_reg190_done;
  wire par_done_reg191_in;
  wire par_done_reg191_write_en;
  wire par_done_reg191_clk;
  wire par_done_reg191_out;
  wire par_done_reg191_done;
  wire par_done_reg192_in;
  wire par_done_reg192_write_en;
  wire par_done_reg192_clk;
  wire par_done_reg192_out;
  wire par_done_reg192_done;
  wire par_done_reg193_in;
  wire par_done_reg193_write_en;
  wire par_done_reg193_clk;
  wire par_done_reg193_out;
  wire par_done_reg193_done;
  wire par_done_reg194_in;
  wire par_done_reg194_write_en;
  wire par_done_reg194_clk;
  wire par_done_reg194_out;
  wire par_done_reg194_done;
  wire par_done_reg195_in;
  wire par_done_reg195_write_en;
  wire par_done_reg195_clk;
  wire par_done_reg195_out;
  wire par_done_reg195_done;
  wire par_done_reg196_in;
  wire par_done_reg196_write_en;
  wire par_done_reg196_clk;
  wire par_done_reg196_out;
  wire par_done_reg196_done;
  wire par_done_reg197_in;
  wire par_done_reg197_write_en;
  wire par_done_reg197_clk;
  wire par_done_reg197_out;
  wire par_done_reg197_done;
  wire par_done_reg198_in;
  wire par_done_reg198_write_en;
  wire par_done_reg198_clk;
  wire par_done_reg198_out;
  wire par_done_reg198_done;
  wire par_done_reg199_in;
  wire par_done_reg199_write_en;
  wire par_done_reg199_clk;
  wire par_done_reg199_out;
  wire par_done_reg199_done;
  wire par_done_reg200_in;
  wire par_done_reg200_write_en;
  wire par_done_reg200_clk;
  wire par_done_reg200_out;
  wire par_done_reg200_done;
  wire par_done_reg201_in;
  wire par_done_reg201_write_en;
  wire par_done_reg201_clk;
  wire par_done_reg201_out;
  wire par_done_reg201_done;
  wire par_done_reg202_in;
  wire par_done_reg202_write_en;
  wire par_done_reg202_clk;
  wire par_done_reg202_out;
  wire par_done_reg202_done;
  wire par_done_reg203_in;
  wire par_done_reg203_write_en;
  wire par_done_reg203_clk;
  wire par_done_reg203_out;
  wire par_done_reg203_done;
  wire par_done_reg204_in;
  wire par_done_reg204_write_en;
  wire par_done_reg204_clk;
  wire par_done_reg204_out;
  wire par_done_reg204_done;
  wire par_reset13_in;
  wire par_reset13_write_en;
  wire par_reset13_clk;
  wire par_reset13_out;
  wire par_reset13_done;
  wire par_done_reg205_in;
  wire par_done_reg205_write_en;
  wire par_done_reg205_clk;
  wire par_done_reg205_out;
  wire par_done_reg205_done;
  wire par_done_reg206_in;
  wire par_done_reg206_write_en;
  wire par_done_reg206_clk;
  wire par_done_reg206_out;
  wire par_done_reg206_done;
  wire par_done_reg207_in;
  wire par_done_reg207_write_en;
  wire par_done_reg207_clk;
  wire par_done_reg207_out;
  wire par_done_reg207_done;
  wire par_done_reg208_in;
  wire par_done_reg208_write_en;
  wire par_done_reg208_clk;
  wire par_done_reg208_out;
  wire par_done_reg208_done;
  wire par_done_reg209_in;
  wire par_done_reg209_write_en;
  wire par_done_reg209_clk;
  wire par_done_reg209_out;
  wire par_done_reg209_done;
  wire par_done_reg210_in;
  wire par_done_reg210_write_en;
  wire par_done_reg210_clk;
  wire par_done_reg210_out;
  wire par_done_reg210_done;
  wire par_done_reg211_in;
  wire par_done_reg211_write_en;
  wire par_done_reg211_clk;
  wire par_done_reg211_out;
  wire par_done_reg211_done;
  wire par_done_reg212_in;
  wire par_done_reg212_write_en;
  wire par_done_reg212_clk;
  wire par_done_reg212_out;
  wire par_done_reg212_done;
  wire par_done_reg213_in;
  wire par_done_reg213_write_en;
  wire par_done_reg213_clk;
  wire par_done_reg213_out;
  wire par_done_reg213_done;
  wire par_done_reg214_in;
  wire par_done_reg214_write_en;
  wire par_done_reg214_clk;
  wire par_done_reg214_out;
  wire par_done_reg214_done;
  wire par_done_reg215_in;
  wire par_done_reg215_write_en;
  wire par_done_reg215_clk;
  wire par_done_reg215_out;
  wire par_done_reg215_done;
  wire par_done_reg216_in;
  wire par_done_reg216_write_en;
  wire par_done_reg216_clk;
  wire par_done_reg216_out;
  wire par_done_reg216_done;
  wire par_done_reg217_in;
  wire par_done_reg217_write_en;
  wire par_done_reg217_clk;
  wire par_done_reg217_out;
  wire par_done_reg217_done;
  wire par_done_reg218_in;
  wire par_done_reg218_write_en;
  wire par_done_reg218_clk;
  wire par_done_reg218_out;
  wire par_done_reg218_done;
  wire par_done_reg219_in;
  wire par_done_reg219_write_en;
  wire par_done_reg219_clk;
  wire par_done_reg219_out;
  wire par_done_reg219_done;
  wire par_done_reg220_in;
  wire par_done_reg220_write_en;
  wire par_done_reg220_clk;
  wire par_done_reg220_out;
  wire par_done_reg220_done;
  wire par_done_reg221_in;
  wire par_done_reg221_write_en;
  wire par_done_reg221_clk;
  wire par_done_reg221_out;
  wire par_done_reg221_done;
  wire par_done_reg222_in;
  wire par_done_reg222_write_en;
  wire par_done_reg222_clk;
  wire par_done_reg222_out;
  wire par_done_reg222_done;
  wire par_done_reg223_in;
  wire par_done_reg223_write_en;
  wire par_done_reg223_clk;
  wire par_done_reg223_out;
  wire par_done_reg223_done;
  wire par_done_reg224_in;
  wire par_done_reg224_write_en;
  wire par_done_reg224_clk;
  wire par_done_reg224_out;
  wire par_done_reg224_done;
  wire par_done_reg225_in;
  wire par_done_reg225_write_en;
  wire par_done_reg225_clk;
  wire par_done_reg225_out;
  wire par_done_reg225_done;
  wire par_done_reg226_in;
  wire par_done_reg226_write_en;
  wire par_done_reg226_clk;
  wire par_done_reg226_out;
  wire par_done_reg226_done;
  wire par_done_reg227_in;
  wire par_done_reg227_write_en;
  wire par_done_reg227_clk;
  wire par_done_reg227_out;
  wire par_done_reg227_done;
  wire par_done_reg228_in;
  wire par_done_reg228_write_en;
  wire par_done_reg228_clk;
  wire par_done_reg228_out;
  wire par_done_reg228_done;
  wire par_done_reg229_in;
  wire par_done_reg229_write_en;
  wire par_done_reg229_clk;
  wire par_done_reg229_out;
  wire par_done_reg229_done;
  wire par_done_reg230_in;
  wire par_done_reg230_write_en;
  wire par_done_reg230_clk;
  wire par_done_reg230_out;
  wire par_done_reg230_done;
  wire par_done_reg231_in;
  wire par_done_reg231_write_en;
  wire par_done_reg231_clk;
  wire par_done_reg231_out;
  wire par_done_reg231_done;
  wire par_done_reg232_in;
  wire par_done_reg232_write_en;
  wire par_done_reg232_clk;
  wire par_done_reg232_out;
  wire par_done_reg232_done;
  wire par_done_reg233_in;
  wire par_done_reg233_write_en;
  wire par_done_reg233_clk;
  wire par_done_reg233_out;
  wire par_done_reg233_done;
  wire par_done_reg234_in;
  wire par_done_reg234_write_en;
  wire par_done_reg234_clk;
  wire par_done_reg234_out;
  wire par_done_reg234_done;
  wire par_done_reg235_in;
  wire par_done_reg235_write_en;
  wire par_done_reg235_clk;
  wire par_done_reg235_out;
  wire par_done_reg235_done;
  wire par_done_reg236_in;
  wire par_done_reg236_write_en;
  wire par_done_reg236_clk;
  wire par_done_reg236_out;
  wire par_done_reg236_done;
  wire par_done_reg237_in;
  wire par_done_reg237_write_en;
  wire par_done_reg237_clk;
  wire par_done_reg237_out;
  wire par_done_reg237_done;
  wire par_done_reg238_in;
  wire par_done_reg238_write_en;
  wire par_done_reg238_clk;
  wire par_done_reg238_out;
  wire par_done_reg238_done;
  wire par_done_reg239_in;
  wire par_done_reg239_write_en;
  wire par_done_reg239_clk;
  wire par_done_reg239_out;
  wire par_done_reg239_done;
  wire par_reset14_in;
  wire par_reset14_write_en;
  wire par_reset14_clk;
  wire par_reset14_out;
  wire par_reset14_done;
  wire par_done_reg240_in;
  wire par_done_reg240_write_en;
  wire par_done_reg240_clk;
  wire par_done_reg240_out;
  wire par_done_reg240_done;
  wire par_done_reg241_in;
  wire par_done_reg241_write_en;
  wire par_done_reg241_clk;
  wire par_done_reg241_out;
  wire par_done_reg241_done;
  wire par_done_reg242_in;
  wire par_done_reg242_write_en;
  wire par_done_reg242_clk;
  wire par_done_reg242_out;
  wire par_done_reg242_done;
  wire par_done_reg243_in;
  wire par_done_reg243_write_en;
  wire par_done_reg243_clk;
  wire par_done_reg243_out;
  wire par_done_reg243_done;
  wire par_done_reg244_in;
  wire par_done_reg244_write_en;
  wire par_done_reg244_clk;
  wire par_done_reg244_out;
  wire par_done_reg244_done;
  wire par_done_reg245_in;
  wire par_done_reg245_write_en;
  wire par_done_reg245_clk;
  wire par_done_reg245_out;
  wire par_done_reg245_done;
  wire par_done_reg246_in;
  wire par_done_reg246_write_en;
  wire par_done_reg246_clk;
  wire par_done_reg246_out;
  wire par_done_reg246_done;
  wire par_done_reg247_in;
  wire par_done_reg247_write_en;
  wire par_done_reg247_clk;
  wire par_done_reg247_out;
  wire par_done_reg247_done;
  wire par_done_reg248_in;
  wire par_done_reg248_write_en;
  wire par_done_reg248_clk;
  wire par_done_reg248_out;
  wire par_done_reg248_done;
  wire par_done_reg249_in;
  wire par_done_reg249_write_en;
  wire par_done_reg249_clk;
  wire par_done_reg249_out;
  wire par_done_reg249_done;
  wire par_done_reg250_in;
  wire par_done_reg250_write_en;
  wire par_done_reg250_clk;
  wire par_done_reg250_out;
  wire par_done_reg250_done;
  wire par_done_reg251_in;
  wire par_done_reg251_write_en;
  wire par_done_reg251_clk;
  wire par_done_reg251_out;
  wire par_done_reg251_done;
  wire par_done_reg252_in;
  wire par_done_reg252_write_en;
  wire par_done_reg252_clk;
  wire par_done_reg252_out;
  wire par_done_reg252_done;
  wire par_done_reg253_in;
  wire par_done_reg253_write_en;
  wire par_done_reg253_clk;
  wire par_done_reg253_out;
  wire par_done_reg253_done;
  wire par_done_reg254_in;
  wire par_done_reg254_write_en;
  wire par_done_reg254_clk;
  wire par_done_reg254_out;
  wire par_done_reg254_done;
  wire par_done_reg255_in;
  wire par_done_reg255_write_en;
  wire par_done_reg255_clk;
  wire par_done_reg255_out;
  wire par_done_reg255_done;
  wire par_done_reg256_in;
  wire par_done_reg256_write_en;
  wire par_done_reg256_clk;
  wire par_done_reg256_out;
  wire par_done_reg256_done;
  wire par_done_reg257_in;
  wire par_done_reg257_write_en;
  wire par_done_reg257_clk;
  wire par_done_reg257_out;
  wire par_done_reg257_done;
  wire par_done_reg258_in;
  wire par_done_reg258_write_en;
  wire par_done_reg258_clk;
  wire par_done_reg258_out;
  wire par_done_reg258_done;
  wire par_done_reg259_in;
  wire par_done_reg259_write_en;
  wire par_done_reg259_clk;
  wire par_done_reg259_out;
  wire par_done_reg259_done;
  wire par_done_reg260_in;
  wire par_done_reg260_write_en;
  wire par_done_reg260_clk;
  wire par_done_reg260_out;
  wire par_done_reg260_done;
  wire par_done_reg261_in;
  wire par_done_reg261_write_en;
  wire par_done_reg261_clk;
  wire par_done_reg261_out;
  wire par_done_reg261_done;
  wire par_done_reg262_in;
  wire par_done_reg262_write_en;
  wire par_done_reg262_clk;
  wire par_done_reg262_out;
  wire par_done_reg262_done;
  wire par_done_reg263_in;
  wire par_done_reg263_write_en;
  wire par_done_reg263_clk;
  wire par_done_reg263_out;
  wire par_done_reg263_done;
  wire par_done_reg264_in;
  wire par_done_reg264_write_en;
  wire par_done_reg264_clk;
  wire par_done_reg264_out;
  wire par_done_reg264_done;
  wire par_done_reg265_in;
  wire par_done_reg265_write_en;
  wire par_done_reg265_clk;
  wire par_done_reg265_out;
  wire par_done_reg265_done;
  wire par_done_reg266_in;
  wire par_done_reg266_write_en;
  wire par_done_reg266_clk;
  wire par_done_reg266_out;
  wire par_done_reg266_done;
  wire par_done_reg267_in;
  wire par_done_reg267_write_en;
  wire par_done_reg267_clk;
  wire par_done_reg267_out;
  wire par_done_reg267_done;
  wire par_done_reg268_in;
  wire par_done_reg268_write_en;
  wire par_done_reg268_clk;
  wire par_done_reg268_out;
  wire par_done_reg268_done;
  wire par_done_reg269_in;
  wire par_done_reg269_write_en;
  wire par_done_reg269_clk;
  wire par_done_reg269_out;
  wire par_done_reg269_done;
  wire par_done_reg270_in;
  wire par_done_reg270_write_en;
  wire par_done_reg270_clk;
  wire par_done_reg270_out;
  wire par_done_reg270_done;
  wire par_done_reg271_in;
  wire par_done_reg271_write_en;
  wire par_done_reg271_clk;
  wire par_done_reg271_out;
  wire par_done_reg271_done;
  wire par_done_reg272_in;
  wire par_done_reg272_write_en;
  wire par_done_reg272_clk;
  wire par_done_reg272_out;
  wire par_done_reg272_done;
  wire par_done_reg273_in;
  wire par_done_reg273_write_en;
  wire par_done_reg273_clk;
  wire par_done_reg273_out;
  wire par_done_reg273_done;
  wire par_done_reg274_in;
  wire par_done_reg274_write_en;
  wire par_done_reg274_clk;
  wire par_done_reg274_out;
  wire par_done_reg274_done;
  wire par_done_reg275_in;
  wire par_done_reg275_write_en;
  wire par_done_reg275_clk;
  wire par_done_reg275_out;
  wire par_done_reg275_done;
  wire par_done_reg276_in;
  wire par_done_reg276_write_en;
  wire par_done_reg276_clk;
  wire par_done_reg276_out;
  wire par_done_reg276_done;
  wire par_done_reg277_in;
  wire par_done_reg277_write_en;
  wire par_done_reg277_clk;
  wire par_done_reg277_out;
  wire par_done_reg277_done;
  wire par_done_reg278_in;
  wire par_done_reg278_write_en;
  wire par_done_reg278_clk;
  wire par_done_reg278_out;
  wire par_done_reg278_done;
  wire par_done_reg279_in;
  wire par_done_reg279_write_en;
  wire par_done_reg279_clk;
  wire par_done_reg279_out;
  wire par_done_reg279_done;
  wire par_done_reg280_in;
  wire par_done_reg280_write_en;
  wire par_done_reg280_clk;
  wire par_done_reg280_out;
  wire par_done_reg280_done;
  wire par_done_reg281_in;
  wire par_done_reg281_write_en;
  wire par_done_reg281_clk;
  wire par_done_reg281_out;
  wire par_done_reg281_done;
  wire par_done_reg282_in;
  wire par_done_reg282_write_en;
  wire par_done_reg282_clk;
  wire par_done_reg282_out;
  wire par_done_reg282_done;
  wire par_done_reg283_in;
  wire par_done_reg283_write_en;
  wire par_done_reg283_clk;
  wire par_done_reg283_out;
  wire par_done_reg283_done;
  wire par_done_reg284_in;
  wire par_done_reg284_write_en;
  wire par_done_reg284_clk;
  wire par_done_reg284_out;
  wire par_done_reg284_done;
  wire par_done_reg285_in;
  wire par_done_reg285_write_en;
  wire par_done_reg285_clk;
  wire par_done_reg285_out;
  wire par_done_reg285_done;
  wire par_done_reg286_in;
  wire par_done_reg286_write_en;
  wire par_done_reg286_clk;
  wire par_done_reg286_out;
  wire par_done_reg286_done;
  wire par_done_reg287_in;
  wire par_done_reg287_write_en;
  wire par_done_reg287_clk;
  wire par_done_reg287_out;
  wire par_done_reg287_done;
  wire par_done_reg288_in;
  wire par_done_reg288_write_en;
  wire par_done_reg288_clk;
  wire par_done_reg288_out;
  wire par_done_reg288_done;
  wire par_done_reg289_in;
  wire par_done_reg289_write_en;
  wire par_done_reg289_clk;
  wire par_done_reg289_out;
  wire par_done_reg289_done;
  wire par_done_reg290_in;
  wire par_done_reg290_write_en;
  wire par_done_reg290_clk;
  wire par_done_reg290_out;
  wire par_done_reg290_done;
  wire par_done_reg291_in;
  wire par_done_reg291_write_en;
  wire par_done_reg291_clk;
  wire par_done_reg291_out;
  wire par_done_reg291_done;
  wire par_done_reg292_in;
  wire par_done_reg292_write_en;
  wire par_done_reg292_clk;
  wire par_done_reg292_out;
  wire par_done_reg292_done;
  wire par_done_reg293_in;
  wire par_done_reg293_write_en;
  wire par_done_reg293_clk;
  wire par_done_reg293_out;
  wire par_done_reg293_done;
  wire par_done_reg294_in;
  wire par_done_reg294_write_en;
  wire par_done_reg294_clk;
  wire par_done_reg294_out;
  wire par_done_reg294_done;
  wire par_done_reg295_in;
  wire par_done_reg295_write_en;
  wire par_done_reg295_clk;
  wire par_done_reg295_out;
  wire par_done_reg295_done;
  wire par_reset15_in;
  wire par_reset15_write_en;
  wire par_reset15_clk;
  wire par_reset15_out;
  wire par_reset15_done;
  wire par_done_reg296_in;
  wire par_done_reg296_write_en;
  wire par_done_reg296_clk;
  wire par_done_reg296_out;
  wire par_done_reg296_done;
  wire par_done_reg297_in;
  wire par_done_reg297_write_en;
  wire par_done_reg297_clk;
  wire par_done_reg297_out;
  wire par_done_reg297_done;
  wire par_done_reg298_in;
  wire par_done_reg298_write_en;
  wire par_done_reg298_clk;
  wire par_done_reg298_out;
  wire par_done_reg298_done;
  wire par_done_reg299_in;
  wire par_done_reg299_write_en;
  wire par_done_reg299_clk;
  wire par_done_reg299_out;
  wire par_done_reg299_done;
  wire par_done_reg300_in;
  wire par_done_reg300_write_en;
  wire par_done_reg300_clk;
  wire par_done_reg300_out;
  wire par_done_reg300_done;
  wire par_done_reg301_in;
  wire par_done_reg301_write_en;
  wire par_done_reg301_clk;
  wire par_done_reg301_out;
  wire par_done_reg301_done;
  wire par_done_reg302_in;
  wire par_done_reg302_write_en;
  wire par_done_reg302_clk;
  wire par_done_reg302_out;
  wire par_done_reg302_done;
  wire par_done_reg303_in;
  wire par_done_reg303_write_en;
  wire par_done_reg303_clk;
  wire par_done_reg303_out;
  wire par_done_reg303_done;
  wire par_done_reg304_in;
  wire par_done_reg304_write_en;
  wire par_done_reg304_clk;
  wire par_done_reg304_out;
  wire par_done_reg304_done;
  wire par_done_reg305_in;
  wire par_done_reg305_write_en;
  wire par_done_reg305_clk;
  wire par_done_reg305_out;
  wire par_done_reg305_done;
  wire par_done_reg306_in;
  wire par_done_reg306_write_en;
  wire par_done_reg306_clk;
  wire par_done_reg306_out;
  wire par_done_reg306_done;
  wire par_done_reg307_in;
  wire par_done_reg307_write_en;
  wire par_done_reg307_clk;
  wire par_done_reg307_out;
  wire par_done_reg307_done;
  wire par_done_reg308_in;
  wire par_done_reg308_write_en;
  wire par_done_reg308_clk;
  wire par_done_reg308_out;
  wire par_done_reg308_done;
  wire par_done_reg309_in;
  wire par_done_reg309_write_en;
  wire par_done_reg309_clk;
  wire par_done_reg309_out;
  wire par_done_reg309_done;
  wire par_done_reg310_in;
  wire par_done_reg310_write_en;
  wire par_done_reg310_clk;
  wire par_done_reg310_out;
  wire par_done_reg310_done;
  wire par_done_reg311_in;
  wire par_done_reg311_write_en;
  wire par_done_reg311_clk;
  wire par_done_reg311_out;
  wire par_done_reg311_done;
  wire par_done_reg312_in;
  wire par_done_reg312_write_en;
  wire par_done_reg312_clk;
  wire par_done_reg312_out;
  wire par_done_reg312_done;
  wire par_done_reg313_in;
  wire par_done_reg313_write_en;
  wire par_done_reg313_clk;
  wire par_done_reg313_out;
  wire par_done_reg313_done;
  wire par_done_reg314_in;
  wire par_done_reg314_write_en;
  wire par_done_reg314_clk;
  wire par_done_reg314_out;
  wire par_done_reg314_done;
  wire par_done_reg315_in;
  wire par_done_reg315_write_en;
  wire par_done_reg315_clk;
  wire par_done_reg315_out;
  wire par_done_reg315_done;
  wire par_done_reg316_in;
  wire par_done_reg316_write_en;
  wire par_done_reg316_clk;
  wire par_done_reg316_out;
  wire par_done_reg316_done;
  wire par_done_reg317_in;
  wire par_done_reg317_write_en;
  wire par_done_reg317_clk;
  wire par_done_reg317_out;
  wire par_done_reg317_done;
  wire par_done_reg318_in;
  wire par_done_reg318_write_en;
  wire par_done_reg318_clk;
  wire par_done_reg318_out;
  wire par_done_reg318_done;
  wire par_done_reg319_in;
  wire par_done_reg319_write_en;
  wire par_done_reg319_clk;
  wire par_done_reg319_out;
  wire par_done_reg319_done;
  wire par_done_reg320_in;
  wire par_done_reg320_write_en;
  wire par_done_reg320_clk;
  wire par_done_reg320_out;
  wire par_done_reg320_done;
  wire par_done_reg321_in;
  wire par_done_reg321_write_en;
  wire par_done_reg321_clk;
  wire par_done_reg321_out;
  wire par_done_reg321_done;
  wire par_done_reg322_in;
  wire par_done_reg322_write_en;
  wire par_done_reg322_clk;
  wire par_done_reg322_out;
  wire par_done_reg322_done;
  wire par_done_reg323_in;
  wire par_done_reg323_write_en;
  wire par_done_reg323_clk;
  wire par_done_reg323_out;
  wire par_done_reg323_done;
  wire par_done_reg324_in;
  wire par_done_reg324_write_en;
  wire par_done_reg324_clk;
  wire par_done_reg324_out;
  wire par_done_reg324_done;
  wire par_done_reg325_in;
  wire par_done_reg325_write_en;
  wire par_done_reg325_clk;
  wire par_done_reg325_out;
  wire par_done_reg325_done;
  wire par_done_reg326_in;
  wire par_done_reg326_write_en;
  wire par_done_reg326_clk;
  wire par_done_reg326_out;
  wire par_done_reg326_done;
  wire par_done_reg327_in;
  wire par_done_reg327_write_en;
  wire par_done_reg327_clk;
  wire par_done_reg327_out;
  wire par_done_reg327_done;
  wire par_done_reg328_in;
  wire par_done_reg328_write_en;
  wire par_done_reg328_clk;
  wire par_done_reg328_out;
  wire par_done_reg328_done;
  wire par_done_reg329_in;
  wire par_done_reg329_write_en;
  wire par_done_reg329_clk;
  wire par_done_reg329_out;
  wire par_done_reg329_done;
  wire par_done_reg330_in;
  wire par_done_reg330_write_en;
  wire par_done_reg330_clk;
  wire par_done_reg330_out;
  wire par_done_reg330_done;
  wire par_done_reg331_in;
  wire par_done_reg331_write_en;
  wire par_done_reg331_clk;
  wire par_done_reg331_out;
  wire par_done_reg331_done;
  wire par_done_reg332_in;
  wire par_done_reg332_write_en;
  wire par_done_reg332_clk;
  wire par_done_reg332_out;
  wire par_done_reg332_done;
  wire par_done_reg333_in;
  wire par_done_reg333_write_en;
  wire par_done_reg333_clk;
  wire par_done_reg333_out;
  wire par_done_reg333_done;
  wire par_done_reg334_in;
  wire par_done_reg334_write_en;
  wire par_done_reg334_clk;
  wire par_done_reg334_out;
  wire par_done_reg334_done;
  wire par_done_reg335_in;
  wire par_done_reg335_write_en;
  wire par_done_reg335_clk;
  wire par_done_reg335_out;
  wire par_done_reg335_done;
  wire par_done_reg336_in;
  wire par_done_reg336_write_en;
  wire par_done_reg336_clk;
  wire par_done_reg336_out;
  wire par_done_reg336_done;
  wire par_done_reg337_in;
  wire par_done_reg337_write_en;
  wire par_done_reg337_clk;
  wire par_done_reg337_out;
  wire par_done_reg337_done;
  wire par_done_reg338_in;
  wire par_done_reg338_write_en;
  wire par_done_reg338_clk;
  wire par_done_reg338_out;
  wire par_done_reg338_done;
  wire par_done_reg339_in;
  wire par_done_reg339_write_en;
  wire par_done_reg339_clk;
  wire par_done_reg339_out;
  wire par_done_reg339_done;
  wire par_reset16_in;
  wire par_reset16_write_en;
  wire par_reset16_clk;
  wire par_reset16_out;
  wire par_reset16_done;
  wire par_done_reg340_in;
  wire par_done_reg340_write_en;
  wire par_done_reg340_clk;
  wire par_done_reg340_out;
  wire par_done_reg340_done;
  wire par_done_reg341_in;
  wire par_done_reg341_write_en;
  wire par_done_reg341_clk;
  wire par_done_reg341_out;
  wire par_done_reg341_done;
  wire par_done_reg342_in;
  wire par_done_reg342_write_en;
  wire par_done_reg342_clk;
  wire par_done_reg342_out;
  wire par_done_reg342_done;
  wire par_done_reg343_in;
  wire par_done_reg343_write_en;
  wire par_done_reg343_clk;
  wire par_done_reg343_out;
  wire par_done_reg343_done;
  wire par_done_reg344_in;
  wire par_done_reg344_write_en;
  wire par_done_reg344_clk;
  wire par_done_reg344_out;
  wire par_done_reg344_done;
  wire par_done_reg345_in;
  wire par_done_reg345_write_en;
  wire par_done_reg345_clk;
  wire par_done_reg345_out;
  wire par_done_reg345_done;
  wire par_done_reg346_in;
  wire par_done_reg346_write_en;
  wire par_done_reg346_clk;
  wire par_done_reg346_out;
  wire par_done_reg346_done;
  wire par_done_reg347_in;
  wire par_done_reg347_write_en;
  wire par_done_reg347_clk;
  wire par_done_reg347_out;
  wire par_done_reg347_done;
  wire par_done_reg348_in;
  wire par_done_reg348_write_en;
  wire par_done_reg348_clk;
  wire par_done_reg348_out;
  wire par_done_reg348_done;
  wire par_done_reg349_in;
  wire par_done_reg349_write_en;
  wire par_done_reg349_clk;
  wire par_done_reg349_out;
  wire par_done_reg349_done;
  wire par_done_reg350_in;
  wire par_done_reg350_write_en;
  wire par_done_reg350_clk;
  wire par_done_reg350_out;
  wire par_done_reg350_done;
  wire par_done_reg351_in;
  wire par_done_reg351_write_en;
  wire par_done_reg351_clk;
  wire par_done_reg351_out;
  wire par_done_reg351_done;
  wire par_done_reg352_in;
  wire par_done_reg352_write_en;
  wire par_done_reg352_clk;
  wire par_done_reg352_out;
  wire par_done_reg352_done;
  wire par_done_reg353_in;
  wire par_done_reg353_write_en;
  wire par_done_reg353_clk;
  wire par_done_reg353_out;
  wire par_done_reg353_done;
  wire par_done_reg354_in;
  wire par_done_reg354_write_en;
  wire par_done_reg354_clk;
  wire par_done_reg354_out;
  wire par_done_reg354_done;
  wire par_done_reg355_in;
  wire par_done_reg355_write_en;
  wire par_done_reg355_clk;
  wire par_done_reg355_out;
  wire par_done_reg355_done;
  wire par_done_reg356_in;
  wire par_done_reg356_write_en;
  wire par_done_reg356_clk;
  wire par_done_reg356_out;
  wire par_done_reg356_done;
  wire par_done_reg357_in;
  wire par_done_reg357_write_en;
  wire par_done_reg357_clk;
  wire par_done_reg357_out;
  wire par_done_reg357_done;
  wire par_done_reg358_in;
  wire par_done_reg358_write_en;
  wire par_done_reg358_clk;
  wire par_done_reg358_out;
  wire par_done_reg358_done;
  wire par_done_reg359_in;
  wire par_done_reg359_write_en;
  wire par_done_reg359_clk;
  wire par_done_reg359_out;
  wire par_done_reg359_done;
  wire par_done_reg360_in;
  wire par_done_reg360_write_en;
  wire par_done_reg360_clk;
  wire par_done_reg360_out;
  wire par_done_reg360_done;
  wire par_done_reg361_in;
  wire par_done_reg361_write_en;
  wire par_done_reg361_clk;
  wire par_done_reg361_out;
  wire par_done_reg361_done;
  wire par_done_reg362_in;
  wire par_done_reg362_write_en;
  wire par_done_reg362_clk;
  wire par_done_reg362_out;
  wire par_done_reg362_done;
  wire par_done_reg363_in;
  wire par_done_reg363_write_en;
  wire par_done_reg363_clk;
  wire par_done_reg363_out;
  wire par_done_reg363_done;
  wire par_done_reg364_in;
  wire par_done_reg364_write_en;
  wire par_done_reg364_clk;
  wire par_done_reg364_out;
  wire par_done_reg364_done;
  wire par_done_reg365_in;
  wire par_done_reg365_write_en;
  wire par_done_reg365_clk;
  wire par_done_reg365_out;
  wire par_done_reg365_done;
  wire par_done_reg366_in;
  wire par_done_reg366_write_en;
  wire par_done_reg366_clk;
  wire par_done_reg366_out;
  wire par_done_reg366_done;
  wire par_done_reg367_in;
  wire par_done_reg367_write_en;
  wire par_done_reg367_clk;
  wire par_done_reg367_out;
  wire par_done_reg367_done;
  wire par_done_reg368_in;
  wire par_done_reg368_write_en;
  wire par_done_reg368_clk;
  wire par_done_reg368_out;
  wire par_done_reg368_done;
  wire par_done_reg369_in;
  wire par_done_reg369_write_en;
  wire par_done_reg369_clk;
  wire par_done_reg369_out;
  wire par_done_reg369_done;
  wire par_done_reg370_in;
  wire par_done_reg370_write_en;
  wire par_done_reg370_clk;
  wire par_done_reg370_out;
  wire par_done_reg370_done;
  wire par_done_reg371_in;
  wire par_done_reg371_write_en;
  wire par_done_reg371_clk;
  wire par_done_reg371_out;
  wire par_done_reg371_done;
  wire par_done_reg372_in;
  wire par_done_reg372_write_en;
  wire par_done_reg372_clk;
  wire par_done_reg372_out;
  wire par_done_reg372_done;
  wire par_done_reg373_in;
  wire par_done_reg373_write_en;
  wire par_done_reg373_clk;
  wire par_done_reg373_out;
  wire par_done_reg373_done;
  wire par_done_reg374_in;
  wire par_done_reg374_write_en;
  wire par_done_reg374_clk;
  wire par_done_reg374_out;
  wire par_done_reg374_done;
  wire par_done_reg375_in;
  wire par_done_reg375_write_en;
  wire par_done_reg375_clk;
  wire par_done_reg375_out;
  wire par_done_reg375_done;
  wire par_done_reg376_in;
  wire par_done_reg376_write_en;
  wire par_done_reg376_clk;
  wire par_done_reg376_out;
  wire par_done_reg376_done;
  wire par_done_reg377_in;
  wire par_done_reg377_write_en;
  wire par_done_reg377_clk;
  wire par_done_reg377_out;
  wire par_done_reg377_done;
  wire par_done_reg378_in;
  wire par_done_reg378_write_en;
  wire par_done_reg378_clk;
  wire par_done_reg378_out;
  wire par_done_reg378_done;
  wire par_done_reg379_in;
  wire par_done_reg379_write_en;
  wire par_done_reg379_clk;
  wire par_done_reg379_out;
  wire par_done_reg379_done;
  wire par_done_reg380_in;
  wire par_done_reg380_write_en;
  wire par_done_reg380_clk;
  wire par_done_reg380_out;
  wire par_done_reg380_done;
  wire par_done_reg381_in;
  wire par_done_reg381_write_en;
  wire par_done_reg381_clk;
  wire par_done_reg381_out;
  wire par_done_reg381_done;
  wire par_done_reg382_in;
  wire par_done_reg382_write_en;
  wire par_done_reg382_clk;
  wire par_done_reg382_out;
  wire par_done_reg382_done;
  wire par_done_reg383_in;
  wire par_done_reg383_write_en;
  wire par_done_reg383_clk;
  wire par_done_reg383_out;
  wire par_done_reg383_done;
  wire par_done_reg384_in;
  wire par_done_reg384_write_en;
  wire par_done_reg384_clk;
  wire par_done_reg384_out;
  wire par_done_reg384_done;
  wire par_done_reg385_in;
  wire par_done_reg385_write_en;
  wire par_done_reg385_clk;
  wire par_done_reg385_out;
  wire par_done_reg385_done;
  wire par_done_reg386_in;
  wire par_done_reg386_write_en;
  wire par_done_reg386_clk;
  wire par_done_reg386_out;
  wire par_done_reg386_done;
  wire par_done_reg387_in;
  wire par_done_reg387_write_en;
  wire par_done_reg387_clk;
  wire par_done_reg387_out;
  wire par_done_reg387_done;
  wire par_done_reg388_in;
  wire par_done_reg388_write_en;
  wire par_done_reg388_clk;
  wire par_done_reg388_out;
  wire par_done_reg388_done;
  wire par_done_reg389_in;
  wire par_done_reg389_write_en;
  wire par_done_reg389_clk;
  wire par_done_reg389_out;
  wire par_done_reg389_done;
  wire par_done_reg390_in;
  wire par_done_reg390_write_en;
  wire par_done_reg390_clk;
  wire par_done_reg390_out;
  wire par_done_reg390_done;
  wire par_done_reg391_in;
  wire par_done_reg391_write_en;
  wire par_done_reg391_clk;
  wire par_done_reg391_out;
  wire par_done_reg391_done;
  wire par_done_reg392_in;
  wire par_done_reg392_write_en;
  wire par_done_reg392_clk;
  wire par_done_reg392_out;
  wire par_done_reg392_done;
  wire par_done_reg393_in;
  wire par_done_reg393_write_en;
  wire par_done_reg393_clk;
  wire par_done_reg393_out;
  wire par_done_reg393_done;
  wire par_done_reg394_in;
  wire par_done_reg394_write_en;
  wire par_done_reg394_clk;
  wire par_done_reg394_out;
  wire par_done_reg394_done;
  wire par_done_reg395_in;
  wire par_done_reg395_write_en;
  wire par_done_reg395_clk;
  wire par_done_reg395_out;
  wire par_done_reg395_done;
  wire par_done_reg396_in;
  wire par_done_reg396_write_en;
  wire par_done_reg396_clk;
  wire par_done_reg396_out;
  wire par_done_reg396_done;
  wire par_done_reg397_in;
  wire par_done_reg397_write_en;
  wire par_done_reg397_clk;
  wire par_done_reg397_out;
  wire par_done_reg397_done;
  wire par_done_reg398_in;
  wire par_done_reg398_write_en;
  wire par_done_reg398_clk;
  wire par_done_reg398_out;
  wire par_done_reg398_done;
  wire par_done_reg399_in;
  wire par_done_reg399_write_en;
  wire par_done_reg399_clk;
  wire par_done_reg399_out;
  wire par_done_reg399_done;
  wire par_done_reg400_in;
  wire par_done_reg400_write_en;
  wire par_done_reg400_clk;
  wire par_done_reg400_out;
  wire par_done_reg400_done;
  wire par_done_reg401_in;
  wire par_done_reg401_write_en;
  wire par_done_reg401_clk;
  wire par_done_reg401_out;
  wire par_done_reg401_done;
  wire par_done_reg402_in;
  wire par_done_reg402_write_en;
  wire par_done_reg402_clk;
  wire par_done_reg402_out;
  wire par_done_reg402_done;
  wire par_done_reg403_in;
  wire par_done_reg403_write_en;
  wire par_done_reg403_clk;
  wire par_done_reg403_out;
  wire par_done_reg403_done;
  wire par_done_reg404_in;
  wire par_done_reg404_write_en;
  wire par_done_reg404_clk;
  wire par_done_reg404_out;
  wire par_done_reg404_done;
  wire par_done_reg405_in;
  wire par_done_reg405_write_en;
  wire par_done_reg405_clk;
  wire par_done_reg405_out;
  wire par_done_reg405_done;
  wire par_done_reg406_in;
  wire par_done_reg406_write_en;
  wire par_done_reg406_clk;
  wire par_done_reg406_out;
  wire par_done_reg406_done;
  wire par_done_reg407_in;
  wire par_done_reg407_write_en;
  wire par_done_reg407_clk;
  wire par_done_reg407_out;
  wire par_done_reg407_done;
  wire par_done_reg408_in;
  wire par_done_reg408_write_en;
  wire par_done_reg408_clk;
  wire par_done_reg408_out;
  wire par_done_reg408_done;
  wire par_done_reg409_in;
  wire par_done_reg409_write_en;
  wire par_done_reg409_clk;
  wire par_done_reg409_out;
  wire par_done_reg409_done;
  wire par_done_reg410_in;
  wire par_done_reg410_write_en;
  wire par_done_reg410_clk;
  wire par_done_reg410_out;
  wire par_done_reg410_done;
  wire par_done_reg411_in;
  wire par_done_reg411_write_en;
  wire par_done_reg411_clk;
  wire par_done_reg411_out;
  wire par_done_reg411_done;
  wire par_reset17_in;
  wire par_reset17_write_en;
  wire par_reset17_clk;
  wire par_reset17_out;
  wire par_reset17_done;
  wire par_done_reg412_in;
  wire par_done_reg412_write_en;
  wire par_done_reg412_clk;
  wire par_done_reg412_out;
  wire par_done_reg412_done;
  wire par_done_reg413_in;
  wire par_done_reg413_write_en;
  wire par_done_reg413_clk;
  wire par_done_reg413_out;
  wire par_done_reg413_done;
  wire par_done_reg414_in;
  wire par_done_reg414_write_en;
  wire par_done_reg414_clk;
  wire par_done_reg414_out;
  wire par_done_reg414_done;
  wire par_done_reg415_in;
  wire par_done_reg415_write_en;
  wire par_done_reg415_clk;
  wire par_done_reg415_out;
  wire par_done_reg415_done;
  wire par_done_reg416_in;
  wire par_done_reg416_write_en;
  wire par_done_reg416_clk;
  wire par_done_reg416_out;
  wire par_done_reg416_done;
  wire par_done_reg417_in;
  wire par_done_reg417_write_en;
  wire par_done_reg417_clk;
  wire par_done_reg417_out;
  wire par_done_reg417_done;
  wire par_done_reg418_in;
  wire par_done_reg418_write_en;
  wire par_done_reg418_clk;
  wire par_done_reg418_out;
  wire par_done_reg418_done;
  wire par_done_reg419_in;
  wire par_done_reg419_write_en;
  wire par_done_reg419_clk;
  wire par_done_reg419_out;
  wire par_done_reg419_done;
  wire par_done_reg420_in;
  wire par_done_reg420_write_en;
  wire par_done_reg420_clk;
  wire par_done_reg420_out;
  wire par_done_reg420_done;
  wire par_done_reg421_in;
  wire par_done_reg421_write_en;
  wire par_done_reg421_clk;
  wire par_done_reg421_out;
  wire par_done_reg421_done;
  wire par_done_reg422_in;
  wire par_done_reg422_write_en;
  wire par_done_reg422_clk;
  wire par_done_reg422_out;
  wire par_done_reg422_done;
  wire par_done_reg423_in;
  wire par_done_reg423_write_en;
  wire par_done_reg423_clk;
  wire par_done_reg423_out;
  wire par_done_reg423_done;
  wire par_done_reg424_in;
  wire par_done_reg424_write_en;
  wire par_done_reg424_clk;
  wire par_done_reg424_out;
  wire par_done_reg424_done;
  wire par_done_reg425_in;
  wire par_done_reg425_write_en;
  wire par_done_reg425_clk;
  wire par_done_reg425_out;
  wire par_done_reg425_done;
  wire par_done_reg426_in;
  wire par_done_reg426_write_en;
  wire par_done_reg426_clk;
  wire par_done_reg426_out;
  wire par_done_reg426_done;
  wire par_done_reg427_in;
  wire par_done_reg427_write_en;
  wire par_done_reg427_clk;
  wire par_done_reg427_out;
  wire par_done_reg427_done;
  wire par_done_reg428_in;
  wire par_done_reg428_write_en;
  wire par_done_reg428_clk;
  wire par_done_reg428_out;
  wire par_done_reg428_done;
  wire par_done_reg429_in;
  wire par_done_reg429_write_en;
  wire par_done_reg429_clk;
  wire par_done_reg429_out;
  wire par_done_reg429_done;
  wire par_done_reg430_in;
  wire par_done_reg430_write_en;
  wire par_done_reg430_clk;
  wire par_done_reg430_out;
  wire par_done_reg430_done;
  wire par_done_reg431_in;
  wire par_done_reg431_write_en;
  wire par_done_reg431_clk;
  wire par_done_reg431_out;
  wire par_done_reg431_done;
  wire par_done_reg432_in;
  wire par_done_reg432_write_en;
  wire par_done_reg432_clk;
  wire par_done_reg432_out;
  wire par_done_reg432_done;
  wire par_done_reg433_in;
  wire par_done_reg433_write_en;
  wire par_done_reg433_clk;
  wire par_done_reg433_out;
  wire par_done_reg433_done;
  wire par_done_reg434_in;
  wire par_done_reg434_write_en;
  wire par_done_reg434_clk;
  wire par_done_reg434_out;
  wire par_done_reg434_done;
  wire par_done_reg435_in;
  wire par_done_reg435_write_en;
  wire par_done_reg435_clk;
  wire par_done_reg435_out;
  wire par_done_reg435_done;
  wire par_done_reg436_in;
  wire par_done_reg436_write_en;
  wire par_done_reg436_clk;
  wire par_done_reg436_out;
  wire par_done_reg436_done;
  wire par_done_reg437_in;
  wire par_done_reg437_write_en;
  wire par_done_reg437_clk;
  wire par_done_reg437_out;
  wire par_done_reg437_done;
  wire par_done_reg438_in;
  wire par_done_reg438_write_en;
  wire par_done_reg438_clk;
  wire par_done_reg438_out;
  wire par_done_reg438_done;
  wire par_done_reg439_in;
  wire par_done_reg439_write_en;
  wire par_done_reg439_clk;
  wire par_done_reg439_out;
  wire par_done_reg439_done;
  wire par_done_reg440_in;
  wire par_done_reg440_write_en;
  wire par_done_reg440_clk;
  wire par_done_reg440_out;
  wire par_done_reg440_done;
  wire par_done_reg441_in;
  wire par_done_reg441_write_en;
  wire par_done_reg441_clk;
  wire par_done_reg441_out;
  wire par_done_reg441_done;
  wire par_done_reg442_in;
  wire par_done_reg442_write_en;
  wire par_done_reg442_clk;
  wire par_done_reg442_out;
  wire par_done_reg442_done;
  wire par_done_reg443_in;
  wire par_done_reg443_write_en;
  wire par_done_reg443_clk;
  wire par_done_reg443_out;
  wire par_done_reg443_done;
  wire par_done_reg444_in;
  wire par_done_reg444_write_en;
  wire par_done_reg444_clk;
  wire par_done_reg444_out;
  wire par_done_reg444_done;
  wire par_done_reg445_in;
  wire par_done_reg445_write_en;
  wire par_done_reg445_clk;
  wire par_done_reg445_out;
  wire par_done_reg445_done;
  wire par_done_reg446_in;
  wire par_done_reg446_write_en;
  wire par_done_reg446_clk;
  wire par_done_reg446_out;
  wire par_done_reg446_done;
  wire par_done_reg447_in;
  wire par_done_reg447_write_en;
  wire par_done_reg447_clk;
  wire par_done_reg447_out;
  wire par_done_reg447_done;
  wire par_done_reg448_in;
  wire par_done_reg448_write_en;
  wire par_done_reg448_clk;
  wire par_done_reg448_out;
  wire par_done_reg448_done;
  wire par_done_reg449_in;
  wire par_done_reg449_write_en;
  wire par_done_reg449_clk;
  wire par_done_reg449_out;
  wire par_done_reg449_done;
  wire par_done_reg450_in;
  wire par_done_reg450_write_en;
  wire par_done_reg450_clk;
  wire par_done_reg450_out;
  wire par_done_reg450_done;
  wire par_done_reg451_in;
  wire par_done_reg451_write_en;
  wire par_done_reg451_clk;
  wire par_done_reg451_out;
  wire par_done_reg451_done;
  wire par_done_reg452_in;
  wire par_done_reg452_write_en;
  wire par_done_reg452_clk;
  wire par_done_reg452_out;
  wire par_done_reg452_done;
  wire par_done_reg453_in;
  wire par_done_reg453_write_en;
  wire par_done_reg453_clk;
  wire par_done_reg453_out;
  wire par_done_reg453_done;
  wire par_done_reg454_in;
  wire par_done_reg454_write_en;
  wire par_done_reg454_clk;
  wire par_done_reg454_out;
  wire par_done_reg454_done;
  wire par_done_reg455_in;
  wire par_done_reg455_write_en;
  wire par_done_reg455_clk;
  wire par_done_reg455_out;
  wire par_done_reg455_done;
  wire par_done_reg456_in;
  wire par_done_reg456_write_en;
  wire par_done_reg456_clk;
  wire par_done_reg456_out;
  wire par_done_reg456_done;
  wire par_done_reg457_in;
  wire par_done_reg457_write_en;
  wire par_done_reg457_clk;
  wire par_done_reg457_out;
  wire par_done_reg457_done;
  wire par_done_reg458_in;
  wire par_done_reg458_write_en;
  wire par_done_reg458_clk;
  wire par_done_reg458_out;
  wire par_done_reg458_done;
  wire par_done_reg459_in;
  wire par_done_reg459_write_en;
  wire par_done_reg459_clk;
  wire par_done_reg459_out;
  wire par_done_reg459_done;
  wire par_done_reg460_in;
  wire par_done_reg460_write_en;
  wire par_done_reg460_clk;
  wire par_done_reg460_out;
  wire par_done_reg460_done;
  wire par_done_reg461_in;
  wire par_done_reg461_write_en;
  wire par_done_reg461_clk;
  wire par_done_reg461_out;
  wire par_done_reg461_done;
  wire par_reset18_in;
  wire par_reset18_write_en;
  wire par_reset18_clk;
  wire par_reset18_out;
  wire par_reset18_done;
  wire par_done_reg462_in;
  wire par_done_reg462_write_en;
  wire par_done_reg462_clk;
  wire par_done_reg462_out;
  wire par_done_reg462_done;
  wire par_done_reg463_in;
  wire par_done_reg463_write_en;
  wire par_done_reg463_clk;
  wire par_done_reg463_out;
  wire par_done_reg463_done;
  wire par_done_reg464_in;
  wire par_done_reg464_write_en;
  wire par_done_reg464_clk;
  wire par_done_reg464_out;
  wire par_done_reg464_done;
  wire par_done_reg465_in;
  wire par_done_reg465_write_en;
  wire par_done_reg465_clk;
  wire par_done_reg465_out;
  wire par_done_reg465_done;
  wire par_done_reg466_in;
  wire par_done_reg466_write_en;
  wire par_done_reg466_clk;
  wire par_done_reg466_out;
  wire par_done_reg466_done;
  wire par_done_reg467_in;
  wire par_done_reg467_write_en;
  wire par_done_reg467_clk;
  wire par_done_reg467_out;
  wire par_done_reg467_done;
  wire par_done_reg468_in;
  wire par_done_reg468_write_en;
  wire par_done_reg468_clk;
  wire par_done_reg468_out;
  wire par_done_reg468_done;
  wire par_done_reg469_in;
  wire par_done_reg469_write_en;
  wire par_done_reg469_clk;
  wire par_done_reg469_out;
  wire par_done_reg469_done;
  wire par_done_reg470_in;
  wire par_done_reg470_write_en;
  wire par_done_reg470_clk;
  wire par_done_reg470_out;
  wire par_done_reg470_done;
  wire par_done_reg471_in;
  wire par_done_reg471_write_en;
  wire par_done_reg471_clk;
  wire par_done_reg471_out;
  wire par_done_reg471_done;
  wire par_done_reg472_in;
  wire par_done_reg472_write_en;
  wire par_done_reg472_clk;
  wire par_done_reg472_out;
  wire par_done_reg472_done;
  wire par_done_reg473_in;
  wire par_done_reg473_write_en;
  wire par_done_reg473_clk;
  wire par_done_reg473_out;
  wire par_done_reg473_done;
  wire par_done_reg474_in;
  wire par_done_reg474_write_en;
  wire par_done_reg474_clk;
  wire par_done_reg474_out;
  wire par_done_reg474_done;
  wire par_done_reg475_in;
  wire par_done_reg475_write_en;
  wire par_done_reg475_clk;
  wire par_done_reg475_out;
  wire par_done_reg475_done;
  wire par_done_reg476_in;
  wire par_done_reg476_write_en;
  wire par_done_reg476_clk;
  wire par_done_reg476_out;
  wire par_done_reg476_done;
  wire par_done_reg477_in;
  wire par_done_reg477_write_en;
  wire par_done_reg477_clk;
  wire par_done_reg477_out;
  wire par_done_reg477_done;
  wire par_done_reg478_in;
  wire par_done_reg478_write_en;
  wire par_done_reg478_clk;
  wire par_done_reg478_out;
  wire par_done_reg478_done;
  wire par_done_reg479_in;
  wire par_done_reg479_write_en;
  wire par_done_reg479_clk;
  wire par_done_reg479_out;
  wire par_done_reg479_done;
  wire par_done_reg480_in;
  wire par_done_reg480_write_en;
  wire par_done_reg480_clk;
  wire par_done_reg480_out;
  wire par_done_reg480_done;
  wire par_done_reg481_in;
  wire par_done_reg481_write_en;
  wire par_done_reg481_clk;
  wire par_done_reg481_out;
  wire par_done_reg481_done;
  wire par_done_reg482_in;
  wire par_done_reg482_write_en;
  wire par_done_reg482_clk;
  wire par_done_reg482_out;
  wire par_done_reg482_done;
  wire par_done_reg483_in;
  wire par_done_reg483_write_en;
  wire par_done_reg483_clk;
  wire par_done_reg483_out;
  wire par_done_reg483_done;
  wire par_done_reg484_in;
  wire par_done_reg484_write_en;
  wire par_done_reg484_clk;
  wire par_done_reg484_out;
  wire par_done_reg484_done;
  wire par_done_reg485_in;
  wire par_done_reg485_write_en;
  wire par_done_reg485_clk;
  wire par_done_reg485_out;
  wire par_done_reg485_done;
  wire par_done_reg486_in;
  wire par_done_reg486_write_en;
  wire par_done_reg486_clk;
  wire par_done_reg486_out;
  wire par_done_reg486_done;
  wire par_done_reg487_in;
  wire par_done_reg487_write_en;
  wire par_done_reg487_clk;
  wire par_done_reg487_out;
  wire par_done_reg487_done;
  wire par_done_reg488_in;
  wire par_done_reg488_write_en;
  wire par_done_reg488_clk;
  wire par_done_reg488_out;
  wire par_done_reg488_done;
  wire par_done_reg489_in;
  wire par_done_reg489_write_en;
  wire par_done_reg489_clk;
  wire par_done_reg489_out;
  wire par_done_reg489_done;
  wire par_done_reg490_in;
  wire par_done_reg490_write_en;
  wire par_done_reg490_clk;
  wire par_done_reg490_out;
  wire par_done_reg490_done;
  wire par_done_reg491_in;
  wire par_done_reg491_write_en;
  wire par_done_reg491_clk;
  wire par_done_reg491_out;
  wire par_done_reg491_done;
  wire par_done_reg492_in;
  wire par_done_reg492_write_en;
  wire par_done_reg492_clk;
  wire par_done_reg492_out;
  wire par_done_reg492_done;
  wire par_done_reg493_in;
  wire par_done_reg493_write_en;
  wire par_done_reg493_clk;
  wire par_done_reg493_out;
  wire par_done_reg493_done;
  wire par_done_reg494_in;
  wire par_done_reg494_write_en;
  wire par_done_reg494_clk;
  wire par_done_reg494_out;
  wire par_done_reg494_done;
  wire par_done_reg495_in;
  wire par_done_reg495_write_en;
  wire par_done_reg495_clk;
  wire par_done_reg495_out;
  wire par_done_reg495_done;
  wire par_done_reg496_in;
  wire par_done_reg496_write_en;
  wire par_done_reg496_clk;
  wire par_done_reg496_out;
  wire par_done_reg496_done;
  wire par_done_reg497_in;
  wire par_done_reg497_write_en;
  wire par_done_reg497_clk;
  wire par_done_reg497_out;
  wire par_done_reg497_done;
  wire par_done_reg498_in;
  wire par_done_reg498_write_en;
  wire par_done_reg498_clk;
  wire par_done_reg498_out;
  wire par_done_reg498_done;
  wire par_done_reg499_in;
  wire par_done_reg499_write_en;
  wire par_done_reg499_clk;
  wire par_done_reg499_out;
  wire par_done_reg499_done;
  wire par_done_reg500_in;
  wire par_done_reg500_write_en;
  wire par_done_reg500_clk;
  wire par_done_reg500_out;
  wire par_done_reg500_done;
  wire par_done_reg501_in;
  wire par_done_reg501_write_en;
  wire par_done_reg501_clk;
  wire par_done_reg501_out;
  wire par_done_reg501_done;
  wire par_done_reg502_in;
  wire par_done_reg502_write_en;
  wire par_done_reg502_clk;
  wire par_done_reg502_out;
  wire par_done_reg502_done;
  wire par_done_reg503_in;
  wire par_done_reg503_write_en;
  wire par_done_reg503_clk;
  wire par_done_reg503_out;
  wire par_done_reg503_done;
  wire par_done_reg504_in;
  wire par_done_reg504_write_en;
  wire par_done_reg504_clk;
  wire par_done_reg504_out;
  wire par_done_reg504_done;
  wire par_done_reg505_in;
  wire par_done_reg505_write_en;
  wire par_done_reg505_clk;
  wire par_done_reg505_out;
  wire par_done_reg505_done;
  wire par_done_reg506_in;
  wire par_done_reg506_write_en;
  wire par_done_reg506_clk;
  wire par_done_reg506_out;
  wire par_done_reg506_done;
  wire par_done_reg507_in;
  wire par_done_reg507_write_en;
  wire par_done_reg507_clk;
  wire par_done_reg507_out;
  wire par_done_reg507_done;
  wire par_done_reg508_in;
  wire par_done_reg508_write_en;
  wire par_done_reg508_clk;
  wire par_done_reg508_out;
  wire par_done_reg508_done;
  wire par_done_reg509_in;
  wire par_done_reg509_write_en;
  wire par_done_reg509_clk;
  wire par_done_reg509_out;
  wire par_done_reg509_done;
  wire par_done_reg510_in;
  wire par_done_reg510_write_en;
  wire par_done_reg510_clk;
  wire par_done_reg510_out;
  wire par_done_reg510_done;
  wire par_done_reg511_in;
  wire par_done_reg511_write_en;
  wire par_done_reg511_clk;
  wire par_done_reg511_out;
  wire par_done_reg511_done;
  wire par_done_reg512_in;
  wire par_done_reg512_write_en;
  wire par_done_reg512_clk;
  wire par_done_reg512_out;
  wire par_done_reg512_done;
  wire par_done_reg513_in;
  wire par_done_reg513_write_en;
  wire par_done_reg513_clk;
  wire par_done_reg513_out;
  wire par_done_reg513_done;
  wire par_done_reg514_in;
  wire par_done_reg514_write_en;
  wire par_done_reg514_clk;
  wire par_done_reg514_out;
  wire par_done_reg514_done;
  wire par_done_reg515_in;
  wire par_done_reg515_write_en;
  wire par_done_reg515_clk;
  wire par_done_reg515_out;
  wire par_done_reg515_done;
  wire par_done_reg516_in;
  wire par_done_reg516_write_en;
  wire par_done_reg516_clk;
  wire par_done_reg516_out;
  wire par_done_reg516_done;
  wire par_done_reg517_in;
  wire par_done_reg517_write_en;
  wire par_done_reg517_clk;
  wire par_done_reg517_out;
  wire par_done_reg517_done;
  wire par_done_reg518_in;
  wire par_done_reg518_write_en;
  wire par_done_reg518_clk;
  wire par_done_reg518_out;
  wire par_done_reg518_done;
  wire par_done_reg519_in;
  wire par_done_reg519_write_en;
  wire par_done_reg519_clk;
  wire par_done_reg519_out;
  wire par_done_reg519_done;
  wire par_done_reg520_in;
  wire par_done_reg520_write_en;
  wire par_done_reg520_clk;
  wire par_done_reg520_out;
  wire par_done_reg520_done;
  wire par_done_reg521_in;
  wire par_done_reg521_write_en;
  wire par_done_reg521_clk;
  wire par_done_reg521_out;
  wire par_done_reg521_done;
  wire par_done_reg522_in;
  wire par_done_reg522_write_en;
  wire par_done_reg522_clk;
  wire par_done_reg522_out;
  wire par_done_reg522_done;
  wire par_done_reg523_in;
  wire par_done_reg523_write_en;
  wire par_done_reg523_clk;
  wire par_done_reg523_out;
  wire par_done_reg523_done;
  wire par_done_reg524_in;
  wire par_done_reg524_write_en;
  wire par_done_reg524_clk;
  wire par_done_reg524_out;
  wire par_done_reg524_done;
  wire par_done_reg525_in;
  wire par_done_reg525_write_en;
  wire par_done_reg525_clk;
  wire par_done_reg525_out;
  wire par_done_reg525_done;
  wire par_done_reg526_in;
  wire par_done_reg526_write_en;
  wire par_done_reg526_clk;
  wire par_done_reg526_out;
  wire par_done_reg526_done;
  wire par_done_reg527_in;
  wire par_done_reg527_write_en;
  wire par_done_reg527_clk;
  wire par_done_reg527_out;
  wire par_done_reg527_done;
  wire par_done_reg528_in;
  wire par_done_reg528_write_en;
  wire par_done_reg528_clk;
  wire par_done_reg528_out;
  wire par_done_reg528_done;
  wire par_done_reg529_in;
  wire par_done_reg529_write_en;
  wire par_done_reg529_clk;
  wire par_done_reg529_out;
  wire par_done_reg529_done;
  wire par_done_reg530_in;
  wire par_done_reg530_write_en;
  wire par_done_reg530_clk;
  wire par_done_reg530_out;
  wire par_done_reg530_done;
  wire par_done_reg531_in;
  wire par_done_reg531_write_en;
  wire par_done_reg531_clk;
  wire par_done_reg531_out;
  wire par_done_reg531_done;
  wire par_done_reg532_in;
  wire par_done_reg532_write_en;
  wire par_done_reg532_clk;
  wire par_done_reg532_out;
  wire par_done_reg532_done;
  wire par_done_reg533_in;
  wire par_done_reg533_write_en;
  wire par_done_reg533_clk;
  wire par_done_reg533_out;
  wire par_done_reg533_done;
  wire par_done_reg534_in;
  wire par_done_reg534_write_en;
  wire par_done_reg534_clk;
  wire par_done_reg534_out;
  wire par_done_reg534_done;
  wire par_done_reg535_in;
  wire par_done_reg535_write_en;
  wire par_done_reg535_clk;
  wire par_done_reg535_out;
  wire par_done_reg535_done;
  wire par_done_reg536_in;
  wire par_done_reg536_write_en;
  wire par_done_reg536_clk;
  wire par_done_reg536_out;
  wire par_done_reg536_done;
  wire par_done_reg537_in;
  wire par_done_reg537_write_en;
  wire par_done_reg537_clk;
  wire par_done_reg537_out;
  wire par_done_reg537_done;
  wire par_done_reg538_in;
  wire par_done_reg538_write_en;
  wire par_done_reg538_clk;
  wire par_done_reg538_out;
  wire par_done_reg538_done;
  wire par_done_reg539_in;
  wire par_done_reg539_write_en;
  wire par_done_reg539_clk;
  wire par_done_reg539_out;
  wire par_done_reg539_done;
  wire par_done_reg540_in;
  wire par_done_reg540_write_en;
  wire par_done_reg540_clk;
  wire par_done_reg540_out;
  wire par_done_reg540_done;
  wire par_done_reg541_in;
  wire par_done_reg541_write_en;
  wire par_done_reg541_clk;
  wire par_done_reg541_out;
  wire par_done_reg541_done;
  wire par_done_reg542_in;
  wire par_done_reg542_write_en;
  wire par_done_reg542_clk;
  wire par_done_reg542_out;
  wire par_done_reg542_done;
  wire par_done_reg543_in;
  wire par_done_reg543_write_en;
  wire par_done_reg543_clk;
  wire par_done_reg543_out;
  wire par_done_reg543_done;
  wire par_done_reg544_in;
  wire par_done_reg544_write_en;
  wire par_done_reg544_clk;
  wire par_done_reg544_out;
  wire par_done_reg544_done;
  wire par_done_reg545_in;
  wire par_done_reg545_write_en;
  wire par_done_reg545_clk;
  wire par_done_reg545_out;
  wire par_done_reg545_done;
  wire par_reset19_in;
  wire par_reset19_write_en;
  wire par_reset19_clk;
  wire par_reset19_out;
  wire par_reset19_done;
  wire par_done_reg546_in;
  wire par_done_reg546_write_en;
  wire par_done_reg546_clk;
  wire par_done_reg546_out;
  wire par_done_reg546_done;
  wire par_done_reg547_in;
  wire par_done_reg547_write_en;
  wire par_done_reg547_clk;
  wire par_done_reg547_out;
  wire par_done_reg547_done;
  wire par_done_reg548_in;
  wire par_done_reg548_write_en;
  wire par_done_reg548_clk;
  wire par_done_reg548_out;
  wire par_done_reg548_done;
  wire par_done_reg549_in;
  wire par_done_reg549_write_en;
  wire par_done_reg549_clk;
  wire par_done_reg549_out;
  wire par_done_reg549_done;
  wire par_done_reg550_in;
  wire par_done_reg550_write_en;
  wire par_done_reg550_clk;
  wire par_done_reg550_out;
  wire par_done_reg550_done;
  wire par_done_reg551_in;
  wire par_done_reg551_write_en;
  wire par_done_reg551_clk;
  wire par_done_reg551_out;
  wire par_done_reg551_done;
  wire par_done_reg552_in;
  wire par_done_reg552_write_en;
  wire par_done_reg552_clk;
  wire par_done_reg552_out;
  wire par_done_reg552_done;
  wire par_done_reg553_in;
  wire par_done_reg553_write_en;
  wire par_done_reg553_clk;
  wire par_done_reg553_out;
  wire par_done_reg553_done;
  wire par_done_reg554_in;
  wire par_done_reg554_write_en;
  wire par_done_reg554_clk;
  wire par_done_reg554_out;
  wire par_done_reg554_done;
  wire par_done_reg555_in;
  wire par_done_reg555_write_en;
  wire par_done_reg555_clk;
  wire par_done_reg555_out;
  wire par_done_reg555_done;
  wire par_done_reg556_in;
  wire par_done_reg556_write_en;
  wire par_done_reg556_clk;
  wire par_done_reg556_out;
  wire par_done_reg556_done;
  wire par_done_reg557_in;
  wire par_done_reg557_write_en;
  wire par_done_reg557_clk;
  wire par_done_reg557_out;
  wire par_done_reg557_done;
  wire par_done_reg558_in;
  wire par_done_reg558_write_en;
  wire par_done_reg558_clk;
  wire par_done_reg558_out;
  wire par_done_reg558_done;
  wire par_done_reg559_in;
  wire par_done_reg559_write_en;
  wire par_done_reg559_clk;
  wire par_done_reg559_out;
  wire par_done_reg559_done;
  wire par_done_reg560_in;
  wire par_done_reg560_write_en;
  wire par_done_reg560_clk;
  wire par_done_reg560_out;
  wire par_done_reg560_done;
  wire par_done_reg561_in;
  wire par_done_reg561_write_en;
  wire par_done_reg561_clk;
  wire par_done_reg561_out;
  wire par_done_reg561_done;
  wire par_done_reg562_in;
  wire par_done_reg562_write_en;
  wire par_done_reg562_clk;
  wire par_done_reg562_out;
  wire par_done_reg562_done;
  wire par_done_reg563_in;
  wire par_done_reg563_write_en;
  wire par_done_reg563_clk;
  wire par_done_reg563_out;
  wire par_done_reg563_done;
  wire par_done_reg564_in;
  wire par_done_reg564_write_en;
  wire par_done_reg564_clk;
  wire par_done_reg564_out;
  wire par_done_reg564_done;
  wire par_done_reg565_in;
  wire par_done_reg565_write_en;
  wire par_done_reg565_clk;
  wire par_done_reg565_out;
  wire par_done_reg565_done;
  wire par_done_reg566_in;
  wire par_done_reg566_write_en;
  wire par_done_reg566_clk;
  wire par_done_reg566_out;
  wire par_done_reg566_done;
  wire par_done_reg567_in;
  wire par_done_reg567_write_en;
  wire par_done_reg567_clk;
  wire par_done_reg567_out;
  wire par_done_reg567_done;
  wire par_done_reg568_in;
  wire par_done_reg568_write_en;
  wire par_done_reg568_clk;
  wire par_done_reg568_out;
  wire par_done_reg568_done;
  wire par_done_reg569_in;
  wire par_done_reg569_write_en;
  wire par_done_reg569_clk;
  wire par_done_reg569_out;
  wire par_done_reg569_done;
  wire par_done_reg570_in;
  wire par_done_reg570_write_en;
  wire par_done_reg570_clk;
  wire par_done_reg570_out;
  wire par_done_reg570_done;
  wire par_done_reg571_in;
  wire par_done_reg571_write_en;
  wire par_done_reg571_clk;
  wire par_done_reg571_out;
  wire par_done_reg571_done;
  wire par_done_reg572_in;
  wire par_done_reg572_write_en;
  wire par_done_reg572_clk;
  wire par_done_reg572_out;
  wire par_done_reg572_done;
  wire par_done_reg573_in;
  wire par_done_reg573_write_en;
  wire par_done_reg573_clk;
  wire par_done_reg573_out;
  wire par_done_reg573_done;
  wire par_done_reg574_in;
  wire par_done_reg574_write_en;
  wire par_done_reg574_clk;
  wire par_done_reg574_out;
  wire par_done_reg574_done;
  wire par_done_reg575_in;
  wire par_done_reg575_write_en;
  wire par_done_reg575_clk;
  wire par_done_reg575_out;
  wire par_done_reg575_done;
  wire par_done_reg576_in;
  wire par_done_reg576_write_en;
  wire par_done_reg576_clk;
  wire par_done_reg576_out;
  wire par_done_reg576_done;
  wire par_done_reg577_in;
  wire par_done_reg577_write_en;
  wire par_done_reg577_clk;
  wire par_done_reg577_out;
  wire par_done_reg577_done;
  wire par_done_reg578_in;
  wire par_done_reg578_write_en;
  wire par_done_reg578_clk;
  wire par_done_reg578_out;
  wire par_done_reg578_done;
  wire par_done_reg579_in;
  wire par_done_reg579_write_en;
  wire par_done_reg579_clk;
  wire par_done_reg579_out;
  wire par_done_reg579_done;
  wire par_done_reg580_in;
  wire par_done_reg580_write_en;
  wire par_done_reg580_clk;
  wire par_done_reg580_out;
  wire par_done_reg580_done;
  wire par_done_reg581_in;
  wire par_done_reg581_write_en;
  wire par_done_reg581_clk;
  wire par_done_reg581_out;
  wire par_done_reg581_done;
  wire par_done_reg582_in;
  wire par_done_reg582_write_en;
  wire par_done_reg582_clk;
  wire par_done_reg582_out;
  wire par_done_reg582_done;
  wire par_done_reg583_in;
  wire par_done_reg583_write_en;
  wire par_done_reg583_clk;
  wire par_done_reg583_out;
  wire par_done_reg583_done;
  wire par_done_reg584_in;
  wire par_done_reg584_write_en;
  wire par_done_reg584_clk;
  wire par_done_reg584_out;
  wire par_done_reg584_done;
  wire par_done_reg585_in;
  wire par_done_reg585_write_en;
  wire par_done_reg585_clk;
  wire par_done_reg585_out;
  wire par_done_reg585_done;
  wire par_done_reg586_in;
  wire par_done_reg586_write_en;
  wire par_done_reg586_clk;
  wire par_done_reg586_out;
  wire par_done_reg586_done;
  wire par_done_reg587_in;
  wire par_done_reg587_write_en;
  wire par_done_reg587_clk;
  wire par_done_reg587_out;
  wire par_done_reg587_done;
  wire par_done_reg588_in;
  wire par_done_reg588_write_en;
  wire par_done_reg588_clk;
  wire par_done_reg588_out;
  wire par_done_reg588_done;
  wire par_done_reg589_in;
  wire par_done_reg589_write_en;
  wire par_done_reg589_clk;
  wire par_done_reg589_out;
  wire par_done_reg589_done;
  wire par_done_reg590_in;
  wire par_done_reg590_write_en;
  wire par_done_reg590_clk;
  wire par_done_reg590_out;
  wire par_done_reg590_done;
  wire par_done_reg591_in;
  wire par_done_reg591_write_en;
  wire par_done_reg591_clk;
  wire par_done_reg591_out;
  wire par_done_reg591_done;
  wire par_done_reg592_in;
  wire par_done_reg592_write_en;
  wire par_done_reg592_clk;
  wire par_done_reg592_out;
  wire par_done_reg592_done;
  wire par_done_reg593_in;
  wire par_done_reg593_write_en;
  wire par_done_reg593_clk;
  wire par_done_reg593_out;
  wire par_done_reg593_done;
  wire par_done_reg594_in;
  wire par_done_reg594_write_en;
  wire par_done_reg594_clk;
  wire par_done_reg594_out;
  wire par_done_reg594_done;
  wire par_done_reg595_in;
  wire par_done_reg595_write_en;
  wire par_done_reg595_clk;
  wire par_done_reg595_out;
  wire par_done_reg595_done;
  wire par_done_reg596_in;
  wire par_done_reg596_write_en;
  wire par_done_reg596_clk;
  wire par_done_reg596_out;
  wire par_done_reg596_done;
  wire par_done_reg597_in;
  wire par_done_reg597_write_en;
  wire par_done_reg597_clk;
  wire par_done_reg597_out;
  wire par_done_reg597_done;
  wire par_done_reg598_in;
  wire par_done_reg598_write_en;
  wire par_done_reg598_clk;
  wire par_done_reg598_out;
  wire par_done_reg598_done;
  wire par_done_reg599_in;
  wire par_done_reg599_write_en;
  wire par_done_reg599_clk;
  wire par_done_reg599_out;
  wire par_done_reg599_done;
  wire par_reset20_in;
  wire par_reset20_write_en;
  wire par_reset20_clk;
  wire par_reset20_out;
  wire par_reset20_done;
  wire par_done_reg600_in;
  wire par_done_reg600_write_en;
  wire par_done_reg600_clk;
  wire par_done_reg600_out;
  wire par_done_reg600_done;
  wire par_done_reg601_in;
  wire par_done_reg601_write_en;
  wire par_done_reg601_clk;
  wire par_done_reg601_out;
  wire par_done_reg601_done;
  wire par_done_reg602_in;
  wire par_done_reg602_write_en;
  wire par_done_reg602_clk;
  wire par_done_reg602_out;
  wire par_done_reg602_done;
  wire par_done_reg603_in;
  wire par_done_reg603_write_en;
  wire par_done_reg603_clk;
  wire par_done_reg603_out;
  wire par_done_reg603_done;
  wire par_done_reg604_in;
  wire par_done_reg604_write_en;
  wire par_done_reg604_clk;
  wire par_done_reg604_out;
  wire par_done_reg604_done;
  wire par_done_reg605_in;
  wire par_done_reg605_write_en;
  wire par_done_reg605_clk;
  wire par_done_reg605_out;
  wire par_done_reg605_done;
  wire par_done_reg606_in;
  wire par_done_reg606_write_en;
  wire par_done_reg606_clk;
  wire par_done_reg606_out;
  wire par_done_reg606_done;
  wire par_done_reg607_in;
  wire par_done_reg607_write_en;
  wire par_done_reg607_clk;
  wire par_done_reg607_out;
  wire par_done_reg607_done;
  wire par_done_reg608_in;
  wire par_done_reg608_write_en;
  wire par_done_reg608_clk;
  wire par_done_reg608_out;
  wire par_done_reg608_done;
  wire par_done_reg609_in;
  wire par_done_reg609_write_en;
  wire par_done_reg609_clk;
  wire par_done_reg609_out;
  wire par_done_reg609_done;
  wire par_done_reg610_in;
  wire par_done_reg610_write_en;
  wire par_done_reg610_clk;
  wire par_done_reg610_out;
  wire par_done_reg610_done;
  wire par_done_reg611_in;
  wire par_done_reg611_write_en;
  wire par_done_reg611_clk;
  wire par_done_reg611_out;
  wire par_done_reg611_done;
  wire par_done_reg612_in;
  wire par_done_reg612_write_en;
  wire par_done_reg612_clk;
  wire par_done_reg612_out;
  wire par_done_reg612_done;
  wire par_done_reg613_in;
  wire par_done_reg613_write_en;
  wire par_done_reg613_clk;
  wire par_done_reg613_out;
  wire par_done_reg613_done;
  wire par_done_reg614_in;
  wire par_done_reg614_write_en;
  wire par_done_reg614_clk;
  wire par_done_reg614_out;
  wire par_done_reg614_done;
  wire par_done_reg615_in;
  wire par_done_reg615_write_en;
  wire par_done_reg615_clk;
  wire par_done_reg615_out;
  wire par_done_reg615_done;
  wire par_done_reg616_in;
  wire par_done_reg616_write_en;
  wire par_done_reg616_clk;
  wire par_done_reg616_out;
  wire par_done_reg616_done;
  wire par_done_reg617_in;
  wire par_done_reg617_write_en;
  wire par_done_reg617_clk;
  wire par_done_reg617_out;
  wire par_done_reg617_done;
  wire par_done_reg618_in;
  wire par_done_reg618_write_en;
  wire par_done_reg618_clk;
  wire par_done_reg618_out;
  wire par_done_reg618_done;
  wire par_done_reg619_in;
  wire par_done_reg619_write_en;
  wire par_done_reg619_clk;
  wire par_done_reg619_out;
  wire par_done_reg619_done;
  wire par_done_reg620_in;
  wire par_done_reg620_write_en;
  wire par_done_reg620_clk;
  wire par_done_reg620_out;
  wire par_done_reg620_done;
  wire par_done_reg621_in;
  wire par_done_reg621_write_en;
  wire par_done_reg621_clk;
  wire par_done_reg621_out;
  wire par_done_reg621_done;
  wire par_done_reg622_in;
  wire par_done_reg622_write_en;
  wire par_done_reg622_clk;
  wire par_done_reg622_out;
  wire par_done_reg622_done;
  wire par_done_reg623_in;
  wire par_done_reg623_write_en;
  wire par_done_reg623_clk;
  wire par_done_reg623_out;
  wire par_done_reg623_done;
  wire par_done_reg624_in;
  wire par_done_reg624_write_en;
  wire par_done_reg624_clk;
  wire par_done_reg624_out;
  wire par_done_reg624_done;
  wire par_done_reg625_in;
  wire par_done_reg625_write_en;
  wire par_done_reg625_clk;
  wire par_done_reg625_out;
  wire par_done_reg625_done;
  wire par_done_reg626_in;
  wire par_done_reg626_write_en;
  wire par_done_reg626_clk;
  wire par_done_reg626_out;
  wire par_done_reg626_done;
  wire par_done_reg627_in;
  wire par_done_reg627_write_en;
  wire par_done_reg627_clk;
  wire par_done_reg627_out;
  wire par_done_reg627_done;
  wire par_done_reg628_in;
  wire par_done_reg628_write_en;
  wire par_done_reg628_clk;
  wire par_done_reg628_out;
  wire par_done_reg628_done;
  wire par_done_reg629_in;
  wire par_done_reg629_write_en;
  wire par_done_reg629_clk;
  wire par_done_reg629_out;
  wire par_done_reg629_done;
  wire par_done_reg630_in;
  wire par_done_reg630_write_en;
  wire par_done_reg630_clk;
  wire par_done_reg630_out;
  wire par_done_reg630_done;
  wire par_done_reg631_in;
  wire par_done_reg631_write_en;
  wire par_done_reg631_clk;
  wire par_done_reg631_out;
  wire par_done_reg631_done;
  wire par_done_reg632_in;
  wire par_done_reg632_write_en;
  wire par_done_reg632_clk;
  wire par_done_reg632_out;
  wire par_done_reg632_done;
  wire par_done_reg633_in;
  wire par_done_reg633_write_en;
  wire par_done_reg633_clk;
  wire par_done_reg633_out;
  wire par_done_reg633_done;
  wire par_done_reg634_in;
  wire par_done_reg634_write_en;
  wire par_done_reg634_clk;
  wire par_done_reg634_out;
  wire par_done_reg634_done;
  wire par_done_reg635_in;
  wire par_done_reg635_write_en;
  wire par_done_reg635_clk;
  wire par_done_reg635_out;
  wire par_done_reg635_done;
  wire par_done_reg636_in;
  wire par_done_reg636_write_en;
  wire par_done_reg636_clk;
  wire par_done_reg636_out;
  wire par_done_reg636_done;
  wire par_done_reg637_in;
  wire par_done_reg637_write_en;
  wire par_done_reg637_clk;
  wire par_done_reg637_out;
  wire par_done_reg637_done;
  wire par_done_reg638_in;
  wire par_done_reg638_write_en;
  wire par_done_reg638_clk;
  wire par_done_reg638_out;
  wire par_done_reg638_done;
  wire par_done_reg639_in;
  wire par_done_reg639_write_en;
  wire par_done_reg639_clk;
  wire par_done_reg639_out;
  wire par_done_reg639_done;
  wire par_done_reg640_in;
  wire par_done_reg640_write_en;
  wire par_done_reg640_clk;
  wire par_done_reg640_out;
  wire par_done_reg640_done;
  wire par_done_reg641_in;
  wire par_done_reg641_write_en;
  wire par_done_reg641_clk;
  wire par_done_reg641_out;
  wire par_done_reg641_done;
  wire par_done_reg642_in;
  wire par_done_reg642_write_en;
  wire par_done_reg642_clk;
  wire par_done_reg642_out;
  wire par_done_reg642_done;
  wire par_done_reg643_in;
  wire par_done_reg643_write_en;
  wire par_done_reg643_clk;
  wire par_done_reg643_out;
  wire par_done_reg643_done;
  wire par_done_reg644_in;
  wire par_done_reg644_write_en;
  wire par_done_reg644_clk;
  wire par_done_reg644_out;
  wire par_done_reg644_done;
  wire par_done_reg645_in;
  wire par_done_reg645_write_en;
  wire par_done_reg645_clk;
  wire par_done_reg645_out;
  wire par_done_reg645_done;
  wire par_done_reg646_in;
  wire par_done_reg646_write_en;
  wire par_done_reg646_clk;
  wire par_done_reg646_out;
  wire par_done_reg646_done;
  wire par_done_reg647_in;
  wire par_done_reg647_write_en;
  wire par_done_reg647_clk;
  wire par_done_reg647_out;
  wire par_done_reg647_done;
  wire par_done_reg648_in;
  wire par_done_reg648_write_en;
  wire par_done_reg648_clk;
  wire par_done_reg648_out;
  wire par_done_reg648_done;
  wire par_done_reg649_in;
  wire par_done_reg649_write_en;
  wire par_done_reg649_clk;
  wire par_done_reg649_out;
  wire par_done_reg649_done;
  wire par_done_reg650_in;
  wire par_done_reg650_write_en;
  wire par_done_reg650_clk;
  wire par_done_reg650_out;
  wire par_done_reg650_done;
  wire par_done_reg651_in;
  wire par_done_reg651_write_en;
  wire par_done_reg651_clk;
  wire par_done_reg651_out;
  wire par_done_reg651_done;
  wire par_done_reg652_in;
  wire par_done_reg652_write_en;
  wire par_done_reg652_clk;
  wire par_done_reg652_out;
  wire par_done_reg652_done;
  wire par_done_reg653_in;
  wire par_done_reg653_write_en;
  wire par_done_reg653_clk;
  wire par_done_reg653_out;
  wire par_done_reg653_done;
  wire par_done_reg654_in;
  wire par_done_reg654_write_en;
  wire par_done_reg654_clk;
  wire par_done_reg654_out;
  wire par_done_reg654_done;
  wire par_done_reg655_in;
  wire par_done_reg655_write_en;
  wire par_done_reg655_clk;
  wire par_done_reg655_out;
  wire par_done_reg655_done;
  wire par_done_reg656_in;
  wire par_done_reg656_write_en;
  wire par_done_reg656_clk;
  wire par_done_reg656_out;
  wire par_done_reg656_done;
  wire par_done_reg657_in;
  wire par_done_reg657_write_en;
  wire par_done_reg657_clk;
  wire par_done_reg657_out;
  wire par_done_reg657_done;
  wire par_done_reg658_in;
  wire par_done_reg658_write_en;
  wire par_done_reg658_clk;
  wire par_done_reg658_out;
  wire par_done_reg658_done;
  wire par_done_reg659_in;
  wire par_done_reg659_write_en;
  wire par_done_reg659_clk;
  wire par_done_reg659_out;
  wire par_done_reg659_done;
  wire par_done_reg660_in;
  wire par_done_reg660_write_en;
  wire par_done_reg660_clk;
  wire par_done_reg660_out;
  wire par_done_reg660_done;
  wire par_done_reg661_in;
  wire par_done_reg661_write_en;
  wire par_done_reg661_clk;
  wire par_done_reg661_out;
  wire par_done_reg661_done;
  wire par_done_reg662_in;
  wire par_done_reg662_write_en;
  wire par_done_reg662_clk;
  wire par_done_reg662_out;
  wire par_done_reg662_done;
  wire par_done_reg663_in;
  wire par_done_reg663_write_en;
  wire par_done_reg663_clk;
  wire par_done_reg663_out;
  wire par_done_reg663_done;
  wire par_done_reg664_in;
  wire par_done_reg664_write_en;
  wire par_done_reg664_clk;
  wire par_done_reg664_out;
  wire par_done_reg664_done;
  wire par_done_reg665_in;
  wire par_done_reg665_write_en;
  wire par_done_reg665_clk;
  wire par_done_reg665_out;
  wire par_done_reg665_done;
  wire par_done_reg666_in;
  wire par_done_reg666_write_en;
  wire par_done_reg666_clk;
  wire par_done_reg666_out;
  wire par_done_reg666_done;
  wire par_done_reg667_in;
  wire par_done_reg667_write_en;
  wire par_done_reg667_clk;
  wire par_done_reg667_out;
  wire par_done_reg667_done;
  wire par_done_reg668_in;
  wire par_done_reg668_write_en;
  wire par_done_reg668_clk;
  wire par_done_reg668_out;
  wire par_done_reg668_done;
  wire par_done_reg669_in;
  wire par_done_reg669_write_en;
  wire par_done_reg669_clk;
  wire par_done_reg669_out;
  wire par_done_reg669_done;
  wire par_done_reg670_in;
  wire par_done_reg670_write_en;
  wire par_done_reg670_clk;
  wire par_done_reg670_out;
  wire par_done_reg670_done;
  wire par_done_reg671_in;
  wire par_done_reg671_write_en;
  wire par_done_reg671_clk;
  wire par_done_reg671_out;
  wire par_done_reg671_done;
  wire par_done_reg672_in;
  wire par_done_reg672_write_en;
  wire par_done_reg672_clk;
  wire par_done_reg672_out;
  wire par_done_reg672_done;
  wire par_done_reg673_in;
  wire par_done_reg673_write_en;
  wire par_done_reg673_clk;
  wire par_done_reg673_out;
  wire par_done_reg673_done;
  wire par_done_reg674_in;
  wire par_done_reg674_write_en;
  wire par_done_reg674_clk;
  wire par_done_reg674_out;
  wire par_done_reg674_done;
  wire par_done_reg675_in;
  wire par_done_reg675_write_en;
  wire par_done_reg675_clk;
  wire par_done_reg675_out;
  wire par_done_reg675_done;
  wire par_done_reg676_in;
  wire par_done_reg676_write_en;
  wire par_done_reg676_clk;
  wire par_done_reg676_out;
  wire par_done_reg676_done;
  wire par_done_reg677_in;
  wire par_done_reg677_write_en;
  wire par_done_reg677_clk;
  wire par_done_reg677_out;
  wire par_done_reg677_done;
  wire par_done_reg678_in;
  wire par_done_reg678_write_en;
  wire par_done_reg678_clk;
  wire par_done_reg678_out;
  wire par_done_reg678_done;
  wire par_done_reg679_in;
  wire par_done_reg679_write_en;
  wire par_done_reg679_clk;
  wire par_done_reg679_out;
  wire par_done_reg679_done;
  wire par_done_reg680_in;
  wire par_done_reg680_write_en;
  wire par_done_reg680_clk;
  wire par_done_reg680_out;
  wire par_done_reg680_done;
  wire par_done_reg681_in;
  wire par_done_reg681_write_en;
  wire par_done_reg681_clk;
  wire par_done_reg681_out;
  wire par_done_reg681_done;
  wire par_done_reg682_in;
  wire par_done_reg682_write_en;
  wire par_done_reg682_clk;
  wire par_done_reg682_out;
  wire par_done_reg682_done;
  wire par_done_reg683_in;
  wire par_done_reg683_write_en;
  wire par_done_reg683_clk;
  wire par_done_reg683_out;
  wire par_done_reg683_done;
  wire par_done_reg684_in;
  wire par_done_reg684_write_en;
  wire par_done_reg684_clk;
  wire par_done_reg684_out;
  wire par_done_reg684_done;
  wire par_done_reg685_in;
  wire par_done_reg685_write_en;
  wire par_done_reg685_clk;
  wire par_done_reg685_out;
  wire par_done_reg685_done;
  wire par_done_reg686_in;
  wire par_done_reg686_write_en;
  wire par_done_reg686_clk;
  wire par_done_reg686_out;
  wire par_done_reg686_done;
  wire par_done_reg687_in;
  wire par_done_reg687_write_en;
  wire par_done_reg687_clk;
  wire par_done_reg687_out;
  wire par_done_reg687_done;
  wire par_done_reg688_in;
  wire par_done_reg688_write_en;
  wire par_done_reg688_clk;
  wire par_done_reg688_out;
  wire par_done_reg688_done;
  wire par_done_reg689_in;
  wire par_done_reg689_write_en;
  wire par_done_reg689_clk;
  wire par_done_reg689_out;
  wire par_done_reg689_done;
  wire par_done_reg690_in;
  wire par_done_reg690_write_en;
  wire par_done_reg690_clk;
  wire par_done_reg690_out;
  wire par_done_reg690_done;
  wire par_done_reg691_in;
  wire par_done_reg691_write_en;
  wire par_done_reg691_clk;
  wire par_done_reg691_out;
  wire par_done_reg691_done;
  wire par_reset21_in;
  wire par_reset21_write_en;
  wire par_reset21_clk;
  wire par_reset21_out;
  wire par_reset21_done;
  wire par_done_reg692_in;
  wire par_done_reg692_write_en;
  wire par_done_reg692_clk;
  wire par_done_reg692_out;
  wire par_done_reg692_done;
  wire par_done_reg693_in;
  wire par_done_reg693_write_en;
  wire par_done_reg693_clk;
  wire par_done_reg693_out;
  wire par_done_reg693_done;
  wire par_done_reg694_in;
  wire par_done_reg694_write_en;
  wire par_done_reg694_clk;
  wire par_done_reg694_out;
  wire par_done_reg694_done;
  wire par_done_reg695_in;
  wire par_done_reg695_write_en;
  wire par_done_reg695_clk;
  wire par_done_reg695_out;
  wire par_done_reg695_done;
  wire par_done_reg696_in;
  wire par_done_reg696_write_en;
  wire par_done_reg696_clk;
  wire par_done_reg696_out;
  wire par_done_reg696_done;
  wire par_done_reg697_in;
  wire par_done_reg697_write_en;
  wire par_done_reg697_clk;
  wire par_done_reg697_out;
  wire par_done_reg697_done;
  wire par_done_reg698_in;
  wire par_done_reg698_write_en;
  wire par_done_reg698_clk;
  wire par_done_reg698_out;
  wire par_done_reg698_done;
  wire par_done_reg699_in;
  wire par_done_reg699_write_en;
  wire par_done_reg699_clk;
  wire par_done_reg699_out;
  wire par_done_reg699_done;
  wire par_done_reg700_in;
  wire par_done_reg700_write_en;
  wire par_done_reg700_clk;
  wire par_done_reg700_out;
  wire par_done_reg700_done;
  wire par_done_reg701_in;
  wire par_done_reg701_write_en;
  wire par_done_reg701_clk;
  wire par_done_reg701_out;
  wire par_done_reg701_done;
  wire par_done_reg702_in;
  wire par_done_reg702_write_en;
  wire par_done_reg702_clk;
  wire par_done_reg702_out;
  wire par_done_reg702_done;
  wire par_done_reg703_in;
  wire par_done_reg703_write_en;
  wire par_done_reg703_clk;
  wire par_done_reg703_out;
  wire par_done_reg703_done;
  wire par_done_reg704_in;
  wire par_done_reg704_write_en;
  wire par_done_reg704_clk;
  wire par_done_reg704_out;
  wire par_done_reg704_done;
  wire par_done_reg705_in;
  wire par_done_reg705_write_en;
  wire par_done_reg705_clk;
  wire par_done_reg705_out;
  wire par_done_reg705_done;
  wire par_done_reg706_in;
  wire par_done_reg706_write_en;
  wire par_done_reg706_clk;
  wire par_done_reg706_out;
  wire par_done_reg706_done;
  wire par_done_reg707_in;
  wire par_done_reg707_write_en;
  wire par_done_reg707_clk;
  wire par_done_reg707_out;
  wire par_done_reg707_done;
  wire par_done_reg708_in;
  wire par_done_reg708_write_en;
  wire par_done_reg708_clk;
  wire par_done_reg708_out;
  wire par_done_reg708_done;
  wire par_done_reg709_in;
  wire par_done_reg709_write_en;
  wire par_done_reg709_clk;
  wire par_done_reg709_out;
  wire par_done_reg709_done;
  wire par_done_reg710_in;
  wire par_done_reg710_write_en;
  wire par_done_reg710_clk;
  wire par_done_reg710_out;
  wire par_done_reg710_done;
  wire par_done_reg711_in;
  wire par_done_reg711_write_en;
  wire par_done_reg711_clk;
  wire par_done_reg711_out;
  wire par_done_reg711_done;
  wire par_done_reg712_in;
  wire par_done_reg712_write_en;
  wire par_done_reg712_clk;
  wire par_done_reg712_out;
  wire par_done_reg712_done;
  wire par_done_reg713_in;
  wire par_done_reg713_write_en;
  wire par_done_reg713_clk;
  wire par_done_reg713_out;
  wire par_done_reg713_done;
  wire par_done_reg714_in;
  wire par_done_reg714_write_en;
  wire par_done_reg714_clk;
  wire par_done_reg714_out;
  wire par_done_reg714_done;
  wire par_done_reg715_in;
  wire par_done_reg715_write_en;
  wire par_done_reg715_clk;
  wire par_done_reg715_out;
  wire par_done_reg715_done;
  wire par_done_reg716_in;
  wire par_done_reg716_write_en;
  wire par_done_reg716_clk;
  wire par_done_reg716_out;
  wire par_done_reg716_done;
  wire par_done_reg717_in;
  wire par_done_reg717_write_en;
  wire par_done_reg717_clk;
  wire par_done_reg717_out;
  wire par_done_reg717_done;
  wire par_done_reg718_in;
  wire par_done_reg718_write_en;
  wire par_done_reg718_clk;
  wire par_done_reg718_out;
  wire par_done_reg718_done;
  wire par_done_reg719_in;
  wire par_done_reg719_write_en;
  wire par_done_reg719_clk;
  wire par_done_reg719_out;
  wire par_done_reg719_done;
  wire par_done_reg720_in;
  wire par_done_reg720_write_en;
  wire par_done_reg720_clk;
  wire par_done_reg720_out;
  wire par_done_reg720_done;
  wire par_done_reg721_in;
  wire par_done_reg721_write_en;
  wire par_done_reg721_clk;
  wire par_done_reg721_out;
  wire par_done_reg721_done;
  wire par_done_reg722_in;
  wire par_done_reg722_write_en;
  wire par_done_reg722_clk;
  wire par_done_reg722_out;
  wire par_done_reg722_done;
  wire par_done_reg723_in;
  wire par_done_reg723_write_en;
  wire par_done_reg723_clk;
  wire par_done_reg723_out;
  wire par_done_reg723_done;
  wire par_done_reg724_in;
  wire par_done_reg724_write_en;
  wire par_done_reg724_clk;
  wire par_done_reg724_out;
  wire par_done_reg724_done;
  wire par_done_reg725_in;
  wire par_done_reg725_write_en;
  wire par_done_reg725_clk;
  wire par_done_reg725_out;
  wire par_done_reg725_done;
  wire par_done_reg726_in;
  wire par_done_reg726_write_en;
  wire par_done_reg726_clk;
  wire par_done_reg726_out;
  wire par_done_reg726_done;
  wire par_done_reg727_in;
  wire par_done_reg727_write_en;
  wire par_done_reg727_clk;
  wire par_done_reg727_out;
  wire par_done_reg727_done;
  wire par_done_reg728_in;
  wire par_done_reg728_write_en;
  wire par_done_reg728_clk;
  wire par_done_reg728_out;
  wire par_done_reg728_done;
  wire par_done_reg729_in;
  wire par_done_reg729_write_en;
  wire par_done_reg729_clk;
  wire par_done_reg729_out;
  wire par_done_reg729_done;
  wire par_done_reg730_in;
  wire par_done_reg730_write_en;
  wire par_done_reg730_clk;
  wire par_done_reg730_out;
  wire par_done_reg730_done;
  wire par_done_reg731_in;
  wire par_done_reg731_write_en;
  wire par_done_reg731_clk;
  wire par_done_reg731_out;
  wire par_done_reg731_done;
  wire par_done_reg732_in;
  wire par_done_reg732_write_en;
  wire par_done_reg732_clk;
  wire par_done_reg732_out;
  wire par_done_reg732_done;
  wire par_done_reg733_in;
  wire par_done_reg733_write_en;
  wire par_done_reg733_clk;
  wire par_done_reg733_out;
  wire par_done_reg733_done;
  wire par_done_reg734_in;
  wire par_done_reg734_write_en;
  wire par_done_reg734_clk;
  wire par_done_reg734_out;
  wire par_done_reg734_done;
  wire par_done_reg735_in;
  wire par_done_reg735_write_en;
  wire par_done_reg735_clk;
  wire par_done_reg735_out;
  wire par_done_reg735_done;
  wire par_done_reg736_in;
  wire par_done_reg736_write_en;
  wire par_done_reg736_clk;
  wire par_done_reg736_out;
  wire par_done_reg736_done;
  wire par_done_reg737_in;
  wire par_done_reg737_write_en;
  wire par_done_reg737_clk;
  wire par_done_reg737_out;
  wire par_done_reg737_done;
  wire par_done_reg738_in;
  wire par_done_reg738_write_en;
  wire par_done_reg738_clk;
  wire par_done_reg738_out;
  wire par_done_reg738_done;
  wire par_done_reg739_in;
  wire par_done_reg739_write_en;
  wire par_done_reg739_clk;
  wire par_done_reg739_out;
  wire par_done_reg739_done;
  wire par_done_reg740_in;
  wire par_done_reg740_write_en;
  wire par_done_reg740_clk;
  wire par_done_reg740_out;
  wire par_done_reg740_done;
  wire par_done_reg741_in;
  wire par_done_reg741_write_en;
  wire par_done_reg741_clk;
  wire par_done_reg741_out;
  wire par_done_reg741_done;
  wire par_done_reg742_in;
  wire par_done_reg742_write_en;
  wire par_done_reg742_clk;
  wire par_done_reg742_out;
  wire par_done_reg742_done;
  wire par_done_reg743_in;
  wire par_done_reg743_write_en;
  wire par_done_reg743_clk;
  wire par_done_reg743_out;
  wire par_done_reg743_done;
  wire par_done_reg744_in;
  wire par_done_reg744_write_en;
  wire par_done_reg744_clk;
  wire par_done_reg744_out;
  wire par_done_reg744_done;
  wire par_done_reg745_in;
  wire par_done_reg745_write_en;
  wire par_done_reg745_clk;
  wire par_done_reg745_out;
  wire par_done_reg745_done;
  wire par_done_reg746_in;
  wire par_done_reg746_write_en;
  wire par_done_reg746_clk;
  wire par_done_reg746_out;
  wire par_done_reg746_done;
  wire par_done_reg747_in;
  wire par_done_reg747_write_en;
  wire par_done_reg747_clk;
  wire par_done_reg747_out;
  wire par_done_reg747_done;
  wire par_reset22_in;
  wire par_reset22_write_en;
  wire par_reset22_clk;
  wire par_reset22_out;
  wire par_reset22_done;
  wire par_done_reg748_in;
  wire par_done_reg748_write_en;
  wire par_done_reg748_clk;
  wire par_done_reg748_out;
  wire par_done_reg748_done;
  wire par_done_reg749_in;
  wire par_done_reg749_write_en;
  wire par_done_reg749_clk;
  wire par_done_reg749_out;
  wire par_done_reg749_done;
  wire par_done_reg750_in;
  wire par_done_reg750_write_en;
  wire par_done_reg750_clk;
  wire par_done_reg750_out;
  wire par_done_reg750_done;
  wire par_done_reg751_in;
  wire par_done_reg751_write_en;
  wire par_done_reg751_clk;
  wire par_done_reg751_out;
  wire par_done_reg751_done;
  wire par_done_reg752_in;
  wire par_done_reg752_write_en;
  wire par_done_reg752_clk;
  wire par_done_reg752_out;
  wire par_done_reg752_done;
  wire par_done_reg753_in;
  wire par_done_reg753_write_en;
  wire par_done_reg753_clk;
  wire par_done_reg753_out;
  wire par_done_reg753_done;
  wire par_done_reg754_in;
  wire par_done_reg754_write_en;
  wire par_done_reg754_clk;
  wire par_done_reg754_out;
  wire par_done_reg754_done;
  wire par_done_reg755_in;
  wire par_done_reg755_write_en;
  wire par_done_reg755_clk;
  wire par_done_reg755_out;
  wire par_done_reg755_done;
  wire par_done_reg756_in;
  wire par_done_reg756_write_en;
  wire par_done_reg756_clk;
  wire par_done_reg756_out;
  wire par_done_reg756_done;
  wire par_done_reg757_in;
  wire par_done_reg757_write_en;
  wire par_done_reg757_clk;
  wire par_done_reg757_out;
  wire par_done_reg757_done;
  wire par_done_reg758_in;
  wire par_done_reg758_write_en;
  wire par_done_reg758_clk;
  wire par_done_reg758_out;
  wire par_done_reg758_done;
  wire par_done_reg759_in;
  wire par_done_reg759_write_en;
  wire par_done_reg759_clk;
  wire par_done_reg759_out;
  wire par_done_reg759_done;
  wire par_done_reg760_in;
  wire par_done_reg760_write_en;
  wire par_done_reg760_clk;
  wire par_done_reg760_out;
  wire par_done_reg760_done;
  wire par_done_reg761_in;
  wire par_done_reg761_write_en;
  wire par_done_reg761_clk;
  wire par_done_reg761_out;
  wire par_done_reg761_done;
  wire par_done_reg762_in;
  wire par_done_reg762_write_en;
  wire par_done_reg762_clk;
  wire par_done_reg762_out;
  wire par_done_reg762_done;
  wire par_done_reg763_in;
  wire par_done_reg763_write_en;
  wire par_done_reg763_clk;
  wire par_done_reg763_out;
  wire par_done_reg763_done;
  wire par_done_reg764_in;
  wire par_done_reg764_write_en;
  wire par_done_reg764_clk;
  wire par_done_reg764_out;
  wire par_done_reg764_done;
  wire par_done_reg765_in;
  wire par_done_reg765_write_en;
  wire par_done_reg765_clk;
  wire par_done_reg765_out;
  wire par_done_reg765_done;
  wire par_done_reg766_in;
  wire par_done_reg766_write_en;
  wire par_done_reg766_clk;
  wire par_done_reg766_out;
  wire par_done_reg766_done;
  wire par_done_reg767_in;
  wire par_done_reg767_write_en;
  wire par_done_reg767_clk;
  wire par_done_reg767_out;
  wire par_done_reg767_done;
  wire par_done_reg768_in;
  wire par_done_reg768_write_en;
  wire par_done_reg768_clk;
  wire par_done_reg768_out;
  wire par_done_reg768_done;
  wire par_done_reg769_in;
  wire par_done_reg769_write_en;
  wire par_done_reg769_clk;
  wire par_done_reg769_out;
  wire par_done_reg769_done;
  wire par_done_reg770_in;
  wire par_done_reg770_write_en;
  wire par_done_reg770_clk;
  wire par_done_reg770_out;
  wire par_done_reg770_done;
  wire par_done_reg771_in;
  wire par_done_reg771_write_en;
  wire par_done_reg771_clk;
  wire par_done_reg771_out;
  wire par_done_reg771_done;
  wire par_done_reg772_in;
  wire par_done_reg772_write_en;
  wire par_done_reg772_clk;
  wire par_done_reg772_out;
  wire par_done_reg772_done;
  wire par_done_reg773_in;
  wire par_done_reg773_write_en;
  wire par_done_reg773_clk;
  wire par_done_reg773_out;
  wire par_done_reg773_done;
  wire par_done_reg774_in;
  wire par_done_reg774_write_en;
  wire par_done_reg774_clk;
  wire par_done_reg774_out;
  wire par_done_reg774_done;
  wire par_done_reg775_in;
  wire par_done_reg775_write_en;
  wire par_done_reg775_clk;
  wire par_done_reg775_out;
  wire par_done_reg775_done;
  wire par_done_reg776_in;
  wire par_done_reg776_write_en;
  wire par_done_reg776_clk;
  wire par_done_reg776_out;
  wire par_done_reg776_done;
  wire par_done_reg777_in;
  wire par_done_reg777_write_en;
  wire par_done_reg777_clk;
  wire par_done_reg777_out;
  wire par_done_reg777_done;
  wire par_done_reg778_in;
  wire par_done_reg778_write_en;
  wire par_done_reg778_clk;
  wire par_done_reg778_out;
  wire par_done_reg778_done;
  wire par_done_reg779_in;
  wire par_done_reg779_write_en;
  wire par_done_reg779_clk;
  wire par_done_reg779_out;
  wire par_done_reg779_done;
  wire par_done_reg780_in;
  wire par_done_reg780_write_en;
  wire par_done_reg780_clk;
  wire par_done_reg780_out;
  wire par_done_reg780_done;
  wire par_done_reg781_in;
  wire par_done_reg781_write_en;
  wire par_done_reg781_clk;
  wire par_done_reg781_out;
  wire par_done_reg781_done;
  wire par_done_reg782_in;
  wire par_done_reg782_write_en;
  wire par_done_reg782_clk;
  wire par_done_reg782_out;
  wire par_done_reg782_done;
  wire par_done_reg783_in;
  wire par_done_reg783_write_en;
  wire par_done_reg783_clk;
  wire par_done_reg783_out;
  wire par_done_reg783_done;
  wire par_done_reg784_in;
  wire par_done_reg784_write_en;
  wire par_done_reg784_clk;
  wire par_done_reg784_out;
  wire par_done_reg784_done;
  wire par_done_reg785_in;
  wire par_done_reg785_write_en;
  wire par_done_reg785_clk;
  wire par_done_reg785_out;
  wire par_done_reg785_done;
  wire par_done_reg786_in;
  wire par_done_reg786_write_en;
  wire par_done_reg786_clk;
  wire par_done_reg786_out;
  wire par_done_reg786_done;
  wire par_done_reg787_in;
  wire par_done_reg787_write_en;
  wire par_done_reg787_clk;
  wire par_done_reg787_out;
  wire par_done_reg787_done;
  wire par_done_reg788_in;
  wire par_done_reg788_write_en;
  wire par_done_reg788_clk;
  wire par_done_reg788_out;
  wire par_done_reg788_done;
  wire par_done_reg789_in;
  wire par_done_reg789_write_en;
  wire par_done_reg789_clk;
  wire par_done_reg789_out;
  wire par_done_reg789_done;
  wire par_done_reg790_in;
  wire par_done_reg790_write_en;
  wire par_done_reg790_clk;
  wire par_done_reg790_out;
  wire par_done_reg790_done;
  wire par_done_reg791_in;
  wire par_done_reg791_write_en;
  wire par_done_reg791_clk;
  wire par_done_reg791_out;
  wire par_done_reg791_done;
  wire par_done_reg792_in;
  wire par_done_reg792_write_en;
  wire par_done_reg792_clk;
  wire par_done_reg792_out;
  wire par_done_reg792_done;
  wire par_done_reg793_in;
  wire par_done_reg793_write_en;
  wire par_done_reg793_clk;
  wire par_done_reg793_out;
  wire par_done_reg793_done;
  wire par_done_reg794_in;
  wire par_done_reg794_write_en;
  wire par_done_reg794_clk;
  wire par_done_reg794_out;
  wire par_done_reg794_done;
  wire par_done_reg795_in;
  wire par_done_reg795_write_en;
  wire par_done_reg795_clk;
  wire par_done_reg795_out;
  wire par_done_reg795_done;
  wire par_done_reg796_in;
  wire par_done_reg796_write_en;
  wire par_done_reg796_clk;
  wire par_done_reg796_out;
  wire par_done_reg796_done;
  wire par_done_reg797_in;
  wire par_done_reg797_write_en;
  wire par_done_reg797_clk;
  wire par_done_reg797_out;
  wire par_done_reg797_done;
  wire par_done_reg798_in;
  wire par_done_reg798_write_en;
  wire par_done_reg798_clk;
  wire par_done_reg798_out;
  wire par_done_reg798_done;
  wire par_done_reg799_in;
  wire par_done_reg799_write_en;
  wire par_done_reg799_clk;
  wire par_done_reg799_out;
  wire par_done_reg799_done;
  wire par_done_reg800_in;
  wire par_done_reg800_write_en;
  wire par_done_reg800_clk;
  wire par_done_reg800_out;
  wire par_done_reg800_done;
  wire par_done_reg801_in;
  wire par_done_reg801_write_en;
  wire par_done_reg801_clk;
  wire par_done_reg801_out;
  wire par_done_reg801_done;
  wire par_done_reg802_in;
  wire par_done_reg802_write_en;
  wire par_done_reg802_clk;
  wire par_done_reg802_out;
  wire par_done_reg802_done;
  wire par_done_reg803_in;
  wire par_done_reg803_write_en;
  wire par_done_reg803_clk;
  wire par_done_reg803_out;
  wire par_done_reg803_done;
  wire par_done_reg804_in;
  wire par_done_reg804_write_en;
  wire par_done_reg804_clk;
  wire par_done_reg804_out;
  wire par_done_reg804_done;
  wire par_done_reg805_in;
  wire par_done_reg805_write_en;
  wire par_done_reg805_clk;
  wire par_done_reg805_out;
  wire par_done_reg805_done;
  wire par_done_reg806_in;
  wire par_done_reg806_write_en;
  wire par_done_reg806_clk;
  wire par_done_reg806_out;
  wire par_done_reg806_done;
  wire par_done_reg807_in;
  wire par_done_reg807_write_en;
  wire par_done_reg807_clk;
  wire par_done_reg807_out;
  wire par_done_reg807_done;
  wire par_done_reg808_in;
  wire par_done_reg808_write_en;
  wire par_done_reg808_clk;
  wire par_done_reg808_out;
  wire par_done_reg808_done;
  wire par_done_reg809_in;
  wire par_done_reg809_write_en;
  wire par_done_reg809_clk;
  wire par_done_reg809_out;
  wire par_done_reg809_done;
  wire par_done_reg810_in;
  wire par_done_reg810_write_en;
  wire par_done_reg810_clk;
  wire par_done_reg810_out;
  wire par_done_reg810_done;
  wire par_done_reg811_in;
  wire par_done_reg811_write_en;
  wire par_done_reg811_clk;
  wire par_done_reg811_out;
  wire par_done_reg811_done;
  wire par_done_reg812_in;
  wire par_done_reg812_write_en;
  wire par_done_reg812_clk;
  wire par_done_reg812_out;
  wire par_done_reg812_done;
  wire par_done_reg813_in;
  wire par_done_reg813_write_en;
  wire par_done_reg813_clk;
  wire par_done_reg813_out;
  wire par_done_reg813_done;
  wire par_done_reg814_in;
  wire par_done_reg814_write_en;
  wire par_done_reg814_clk;
  wire par_done_reg814_out;
  wire par_done_reg814_done;
  wire par_done_reg815_in;
  wire par_done_reg815_write_en;
  wire par_done_reg815_clk;
  wire par_done_reg815_out;
  wire par_done_reg815_done;
  wire par_done_reg816_in;
  wire par_done_reg816_write_en;
  wire par_done_reg816_clk;
  wire par_done_reg816_out;
  wire par_done_reg816_done;
  wire par_done_reg817_in;
  wire par_done_reg817_write_en;
  wire par_done_reg817_clk;
  wire par_done_reg817_out;
  wire par_done_reg817_done;
  wire par_done_reg818_in;
  wire par_done_reg818_write_en;
  wire par_done_reg818_clk;
  wire par_done_reg818_out;
  wire par_done_reg818_done;
  wire par_done_reg819_in;
  wire par_done_reg819_write_en;
  wire par_done_reg819_clk;
  wire par_done_reg819_out;
  wire par_done_reg819_done;
  wire par_done_reg820_in;
  wire par_done_reg820_write_en;
  wire par_done_reg820_clk;
  wire par_done_reg820_out;
  wire par_done_reg820_done;
  wire par_done_reg821_in;
  wire par_done_reg821_write_en;
  wire par_done_reg821_clk;
  wire par_done_reg821_out;
  wire par_done_reg821_done;
  wire par_done_reg822_in;
  wire par_done_reg822_write_en;
  wire par_done_reg822_clk;
  wire par_done_reg822_out;
  wire par_done_reg822_done;
  wire par_done_reg823_in;
  wire par_done_reg823_write_en;
  wire par_done_reg823_clk;
  wire par_done_reg823_out;
  wire par_done_reg823_done;
  wire par_done_reg824_in;
  wire par_done_reg824_write_en;
  wire par_done_reg824_clk;
  wire par_done_reg824_out;
  wire par_done_reg824_done;
  wire par_done_reg825_in;
  wire par_done_reg825_write_en;
  wire par_done_reg825_clk;
  wire par_done_reg825_out;
  wire par_done_reg825_done;
  wire par_done_reg826_in;
  wire par_done_reg826_write_en;
  wire par_done_reg826_clk;
  wire par_done_reg826_out;
  wire par_done_reg826_done;
  wire par_done_reg827_in;
  wire par_done_reg827_write_en;
  wire par_done_reg827_clk;
  wire par_done_reg827_out;
  wire par_done_reg827_done;
  wire par_done_reg828_in;
  wire par_done_reg828_write_en;
  wire par_done_reg828_clk;
  wire par_done_reg828_out;
  wire par_done_reg828_done;
  wire par_done_reg829_in;
  wire par_done_reg829_write_en;
  wire par_done_reg829_clk;
  wire par_done_reg829_out;
  wire par_done_reg829_done;
  wire par_done_reg830_in;
  wire par_done_reg830_write_en;
  wire par_done_reg830_clk;
  wire par_done_reg830_out;
  wire par_done_reg830_done;
  wire par_done_reg831_in;
  wire par_done_reg831_write_en;
  wire par_done_reg831_clk;
  wire par_done_reg831_out;
  wire par_done_reg831_done;
  wire par_done_reg832_in;
  wire par_done_reg832_write_en;
  wire par_done_reg832_clk;
  wire par_done_reg832_out;
  wire par_done_reg832_done;
  wire par_done_reg833_in;
  wire par_done_reg833_write_en;
  wire par_done_reg833_clk;
  wire par_done_reg833_out;
  wire par_done_reg833_done;
  wire par_done_reg834_in;
  wire par_done_reg834_write_en;
  wire par_done_reg834_clk;
  wire par_done_reg834_out;
  wire par_done_reg834_done;
  wire par_done_reg835_in;
  wire par_done_reg835_write_en;
  wire par_done_reg835_clk;
  wire par_done_reg835_out;
  wire par_done_reg835_done;
  wire par_done_reg836_in;
  wire par_done_reg836_write_en;
  wire par_done_reg836_clk;
  wire par_done_reg836_out;
  wire par_done_reg836_done;
  wire par_done_reg837_in;
  wire par_done_reg837_write_en;
  wire par_done_reg837_clk;
  wire par_done_reg837_out;
  wire par_done_reg837_done;
  wire par_done_reg838_in;
  wire par_done_reg838_write_en;
  wire par_done_reg838_clk;
  wire par_done_reg838_out;
  wire par_done_reg838_done;
  wire par_done_reg839_in;
  wire par_done_reg839_write_en;
  wire par_done_reg839_clk;
  wire par_done_reg839_out;
  wire par_done_reg839_done;
  wire par_done_reg840_in;
  wire par_done_reg840_write_en;
  wire par_done_reg840_clk;
  wire par_done_reg840_out;
  wire par_done_reg840_done;
  wire par_done_reg841_in;
  wire par_done_reg841_write_en;
  wire par_done_reg841_clk;
  wire par_done_reg841_out;
  wire par_done_reg841_done;
  wire par_done_reg842_in;
  wire par_done_reg842_write_en;
  wire par_done_reg842_clk;
  wire par_done_reg842_out;
  wire par_done_reg842_done;
  wire par_done_reg843_in;
  wire par_done_reg843_write_en;
  wire par_done_reg843_clk;
  wire par_done_reg843_out;
  wire par_done_reg843_done;
  wire par_reset23_in;
  wire par_reset23_write_en;
  wire par_reset23_clk;
  wire par_reset23_out;
  wire par_reset23_done;
  wire par_done_reg844_in;
  wire par_done_reg844_write_en;
  wire par_done_reg844_clk;
  wire par_done_reg844_out;
  wire par_done_reg844_done;
  wire par_done_reg845_in;
  wire par_done_reg845_write_en;
  wire par_done_reg845_clk;
  wire par_done_reg845_out;
  wire par_done_reg845_done;
  wire par_done_reg846_in;
  wire par_done_reg846_write_en;
  wire par_done_reg846_clk;
  wire par_done_reg846_out;
  wire par_done_reg846_done;
  wire par_done_reg847_in;
  wire par_done_reg847_write_en;
  wire par_done_reg847_clk;
  wire par_done_reg847_out;
  wire par_done_reg847_done;
  wire par_done_reg848_in;
  wire par_done_reg848_write_en;
  wire par_done_reg848_clk;
  wire par_done_reg848_out;
  wire par_done_reg848_done;
  wire par_done_reg849_in;
  wire par_done_reg849_write_en;
  wire par_done_reg849_clk;
  wire par_done_reg849_out;
  wire par_done_reg849_done;
  wire par_done_reg850_in;
  wire par_done_reg850_write_en;
  wire par_done_reg850_clk;
  wire par_done_reg850_out;
  wire par_done_reg850_done;
  wire par_done_reg851_in;
  wire par_done_reg851_write_en;
  wire par_done_reg851_clk;
  wire par_done_reg851_out;
  wire par_done_reg851_done;
  wire par_done_reg852_in;
  wire par_done_reg852_write_en;
  wire par_done_reg852_clk;
  wire par_done_reg852_out;
  wire par_done_reg852_done;
  wire par_done_reg853_in;
  wire par_done_reg853_write_en;
  wire par_done_reg853_clk;
  wire par_done_reg853_out;
  wire par_done_reg853_done;
  wire par_done_reg854_in;
  wire par_done_reg854_write_en;
  wire par_done_reg854_clk;
  wire par_done_reg854_out;
  wire par_done_reg854_done;
  wire par_done_reg855_in;
  wire par_done_reg855_write_en;
  wire par_done_reg855_clk;
  wire par_done_reg855_out;
  wire par_done_reg855_done;
  wire par_done_reg856_in;
  wire par_done_reg856_write_en;
  wire par_done_reg856_clk;
  wire par_done_reg856_out;
  wire par_done_reg856_done;
  wire par_done_reg857_in;
  wire par_done_reg857_write_en;
  wire par_done_reg857_clk;
  wire par_done_reg857_out;
  wire par_done_reg857_done;
  wire par_done_reg858_in;
  wire par_done_reg858_write_en;
  wire par_done_reg858_clk;
  wire par_done_reg858_out;
  wire par_done_reg858_done;
  wire par_done_reg859_in;
  wire par_done_reg859_write_en;
  wire par_done_reg859_clk;
  wire par_done_reg859_out;
  wire par_done_reg859_done;
  wire par_done_reg860_in;
  wire par_done_reg860_write_en;
  wire par_done_reg860_clk;
  wire par_done_reg860_out;
  wire par_done_reg860_done;
  wire par_done_reg861_in;
  wire par_done_reg861_write_en;
  wire par_done_reg861_clk;
  wire par_done_reg861_out;
  wire par_done_reg861_done;
  wire par_done_reg862_in;
  wire par_done_reg862_write_en;
  wire par_done_reg862_clk;
  wire par_done_reg862_out;
  wire par_done_reg862_done;
  wire par_done_reg863_in;
  wire par_done_reg863_write_en;
  wire par_done_reg863_clk;
  wire par_done_reg863_out;
  wire par_done_reg863_done;
  wire par_done_reg864_in;
  wire par_done_reg864_write_en;
  wire par_done_reg864_clk;
  wire par_done_reg864_out;
  wire par_done_reg864_done;
  wire par_done_reg865_in;
  wire par_done_reg865_write_en;
  wire par_done_reg865_clk;
  wire par_done_reg865_out;
  wire par_done_reg865_done;
  wire par_done_reg866_in;
  wire par_done_reg866_write_en;
  wire par_done_reg866_clk;
  wire par_done_reg866_out;
  wire par_done_reg866_done;
  wire par_done_reg867_in;
  wire par_done_reg867_write_en;
  wire par_done_reg867_clk;
  wire par_done_reg867_out;
  wire par_done_reg867_done;
  wire par_done_reg868_in;
  wire par_done_reg868_write_en;
  wire par_done_reg868_clk;
  wire par_done_reg868_out;
  wire par_done_reg868_done;
  wire par_done_reg869_in;
  wire par_done_reg869_write_en;
  wire par_done_reg869_clk;
  wire par_done_reg869_out;
  wire par_done_reg869_done;
  wire par_done_reg870_in;
  wire par_done_reg870_write_en;
  wire par_done_reg870_clk;
  wire par_done_reg870_out;
  wire par_done_reg870_done;
  wire par_done_reg871_in;
  wire par_done_reg871_write_en;
  wire par_done_reg871_clk;
  wire par_done_reg871_out;
  wire par_done_reg871_done;
  wire par_done_reg872_in;
  wire par_done_reg872_write_en;
  wire par_done_reg872_clk;
  wire par_done_reg872_out;
  wire par_done_reg872_done;
  wire par_done_reg873_in;
  wire par_done_reg873_write_en;
  wire par_done_reg873_clk;
  wire par_done_reg873_out;
  wire par_done_reg873_done;
  wire par_done_reg874_in;
  wire par_done_reg874_write_en;
  wire par_done_reg874_clk;
  wire par_done_reg874_out;
  wire par_done_reg874_done;
  wire par_done_reg875_in;
  wire par_done_reg875_write_en;
  wire par_done_reg875_clk;
  wire par_done_reg875_out;
  wire par_done_reg875_done;
  wire par_done_reg876_in;
  wire par_done_reg876_write_en;
  wire par_done_reg876_clk;
  wire par_done_reg876_out;
  wire par_done_reg876_done;
  wire par_done_reg877_in;
  wire par_done_reg877_write_en;
  wire par_done_reg877_clk;
  wire par_done_reg877_out;
  wire par_done_reg877_done;
  wire par_done_reg878_in;
  wire par_done_reg878_write_en;
  wire par_done_reg878_clk;
  wire par_done_reg878_out;
  wire par_done_reg878_done;
  wire par_done_reg879_in;
  wire par_done_reg879_write_en;
  wire par_done_reg879_clk;
  wire par_done_reg879_out;
  wire par_done_reg879_done;
  wire par_done_reg880_in;
  wire par_done_reg880_write_en;
  wire par_done_reg880_clk;
  wire par_done_reg880_out;
  wire par_done_reg880_done;
  wire par_done_reg881_in;
  wire par_done_reg881_write_en;
  wire par_done_reg881_clk;
  wire par_done_reg881_out;
  wire par_done_reg881_done;
  wire par_done_reg882_in;
  wire par_done_reg882_write_en;
  wire par_done_reg882_clk;
  wire par_done_reg882_out;
  wire par_done_reg882_done;
  wire par_done_reg883_in;
  wire par_done_reg883_write_en;
  wire par_done_reg883_clk;
  wire par_done_reg883_out;
  wire par_done_reg883_done;
  wire par_done_reg884_in;
  wire par_done_reg884_write_en;
  wire par_done_reg884_clk;
  wire par_done_reg884_out;
  wire par_done_reg884_done;
  wire par_done_reg885_in;
  wire par_done_reg885_write_en;
  wire par_done_reg885_clk;
  wire par_done_reg885_out;
  wire par_done_reg885_done;
  wire par_done_reg886_in;
  wire par_done_reg886_write_en;
  wire par_done_reg886_clk;
  wire par_done_reg886_out;
  wire par_done_reg886_done;
  wire par_done_reg887_in;
  wire par_done_reg887_write_en;
  wire par_done_reg887_clk;
  wire par_done_reg887_out;
  wire par_done_reg887_done;
  wire par_done_reg888_in;
  wire par_done_reg888_write_en;
  wire par_done_reg888_clk;
  wire par_done_reg888_out;
  wire par_done_reg888_done;
  wire par_done_reg889_in;
  wire par_done_reg889_write_en;
  wire par_done_reg889_clk;
  wire par_done_reg889_out;
  wire par_done_reg889_done;
  wire par_done_reg890_in;
  wire par_done_reg890_write_en;
  wire par_done_reg890_clk;
  wire par_done_reg890_out;
  wire par_done_reg890_done;
  wire par_done_reg891_in;
  wire par_done_reg891_write_en;
  wire par_done_reg891_clk;
  wire par_done_reg891_out;
  wire par_done_reg891_done;
  wire par_done_reg892_in;
  wire par_done_reg892_write_en;
  wire par_done_reg892_clk;
  wire par_done_reg892_out;
  wire par_done_reg892_done;
  wire par_done_reg893_in;
  wire par_done_reg893_write_en;
  wire par_done_reg893_clk;
  wire par_done_reg893_out;
  wire par_done_reg893_done;
  wire par_done_reg894_in;
  wire par_done_reg894_write_en;
  wire par_done_reg894_clk;
  wire par_done_reg894_out;
  wire par_done_reg894_done;
  wire par_done_reg895_in;
  wire par_done_reg895_write_en;
  wire par_done_reg895_clk;
  wire par_done_reg895_out;
  wire par_done_reg895_done;
  wire par_done_reg896_in;
  wire par_done_reg896_write_en;
  wire par_done_reg896_clk;
  wire par_done_reg896_out;
  wire par_done_reg896_done;
  wire par_done_reg897_in;
  wire par_done_reg897_write_en;
  wire par_done_reg897_clk;
  wire par_done_reg897_out;
  wire par_done_reg897_done;
  wire par_done_reg898_in;
  wire par_done_reg898_write_en;
  wire par_done_reg898_clk;
  wire par_done_reg898_out;
  wire par_done_reg898_done;
  wire par_done_reg899_in;
  wire par_done_reg899_write_en;
  wire par_done_reg899_clk;
  wire par_done_reg899_out;
  wire par_done_reg899_done;
  wire par_reset24_in;
  wire par_reset24_write_en;
  wire par_reset24_clk;
  wire par_reset24_out;
  wire par_reset24_done;
  wire par_done_reg900_in;
  wire par_done_reg900_write_en;
  wire par_done_reg900_clk;
  wire par_done_reg900_out;
  wire par_done_reg900_done;
  wire par_done_reg901_in;
  wire par_done_reg901_write_en;
  wire par_done_reg901_clk;
  wire par_done_reg901_out;
  wire par_done_reg901_done;
  wire par_done_reg902_in;
  wire par_done_reg902_write_en;
  wire par_done_reg902_clk;
  wire par_done_reg902_out;
  wire par_done_reg902_done;
  wire par_done_reg903_in;
  wire par_done_reg903_write_en;
  wire par_done_reg903_clk;
  wire par_done_reg903_out;
  wire par_done_reg903_done;
  wire par_done_reg904_in;
  wire par_done_reg904_write_en;
  wire par_done_reg904_clk;
  wire par_done_reg904_out;
  wire par_done_reg904_done;
  wire par_done_reg905_in;
  wire par_done_reg905_write_en;
  wire par_done_reg905_clk;
  wire par_done_reg905_out;
  wire par_done_reg905_done;
  wire par_done_reg906_in;
  wire par_done_reg906_write_en;
  wire par_done_reg906_clk;
  wire par_done_reg906_out;
  wire par_done_reg906_done;
  wire par_done_reg907_in;
  wire par_done_reg907_write_en;
  wire par_done_reg907_clk;
  wire par_done_reg907_out;
  wire par_done_reg907_done;
  wire par_done_reg908_in;
  wire par_done_reg908_write_en;
  wire par_done_reg908_clk;
  wire par_done_reg908_out;
  wire par_done_reg908_done;
  wire par_done_reg909_in;
  wire par_done_reg909_write_en;
  wire par_done_reg909_clk;
  wire par_done_reg909_out;
  wire par_done_reg909_done;
  wire par_done_reg910_in;
  wire par_done_reg910_write_en;
  wire par_done_reg910_clk;
  wire par_done_reg910_out;
  wire par_done_reg910_done;
  wire par_done_reg911_in;
  wire par_done_reg911_write_en;
  wire par_done_reg911_clk;
  wire par_done_reg911_out;
  wire par_done_reg911_done;
  wire par_done_reg912_in;
  wire par_done_reg912_write_en;
  wire par_done_reg912_clk;
  wire par_done_reg912_out;
  wire par_done_reg912_done;
  wire par_done_reg913_in;
  wire par_done_reg913_write_en;
  wire par_done_reg913_clk;
  wire par_done_reg913_out;
  wire par_done_reg913_done;
  wire par_done_reg914_in;
  wire par_done_reg914_write_en;
  wire par_done_reg914_clk;
  wire par_done_reg914_out;
  wire par_done_reg914_done;
  wire par_done_reg915_in;
  wire par_done_reg915_write_en;
  wire par_done_reg915_clk;
  wire par_done_reg915_out;
  wire par_done_reg915_done;
  wire par_done_reg916_in;
  wire par_done_reg916_write_en;
  wire par_done_reg916_clk;
  wire par_done_reg916_out;
  wire par_done_reg916_done;
  wire par_done_reg917_in;
  wire par_done_reg917_write_en;
  wire par_done_reg917_clk;
  wire par_done_reg917_out;
  wire par_done_reg917_done;
  wire par_done_reg918_in;
  wire par_done_reg918_write_en;
  wire par_done_reg918_clk;
  wire par_done_reg918_out;
  wire par_done_reg918_done;
  wire par_done_reg919_in;
  wire par_done_reg919_write_en;
  wire par_done_reg919_clk;
  wire par_done_reg919_out;
  wire par_done_reg919_done;
  wire par_done_reg920_in;
  wire par_done_reg920_write_en;
  wire par_done_reg920_clk;
  wire par_done_reg920_out;
  wire par_done_reg920_done;
  wire par_done_reg921_in;
  wire par_done_reg921_write_en;
  wire par_done_reg921_clk;
  wire par_done_reg921_out;
  wire par_done_reg921_done;
  wire par_done_reg922_in;
  wire par_done_reg922_write_en;
  wire par_done_reg922_clk;
  wire par_done_reg922_out;
  wire par_done_reg922_done;
  wire par_done_reg923_in;
  wire par_done_reg923_write_en;
  wire par_done_reg923_clk;
  wire par_done_reg923_out;
  wire par_done_reg923_done;
  wire par_done_reg924_in;
  wire par_done_reg924_write_en;
  wire par_done_reg924_clk;
  wire par_done_reg924_out;
  wire par_done_reg924_done;
  wire par_done_reg925_in;
  wire par_done_reg925_write_en;
  wire par_done_reg925_clk;
  wire par_done_reg925_out;
  wire par_done_reg925_done;
  wire par_done_reg926_in;
  wire par_done_reg926_write_en;
  wire par_done_reg926_clk;
  wire par_done_reg926_out;
  wire par_done_reg926_done;
  wire par_done_reg927_in;
  wire par_done_reg927_write_en;
  wire par_done_reg927_clk;
  wire par_done_reg927_out;
  wire par_done_reg927_done;
  wire par_done_reg928_in;
  wire par_done_reg928_write_en;
  wire par_done_reg928_clk;
  wire par_done_reg928_out;
  wire par_done_reg928_done;
  wire par_done_reg929_in;
  wire par_done_reg929_write_en;
  wire par_done_reg929_clk;
  wire par_done_reg929_out;
  wire par_done_reg929_done;
  wire par_done_reg930_in;
  wire par_done_reg930_write_en;
  wire par_done_reg930_clk;
  wire par_done_reg930_out;
  wire par_done_reg930_done;
  wire par_done_reg931_in;
  wire par_done_reg931_write_en;
  wire par_done_reg931_clk;
  wire par_done_reg931_out;
  wire par_done_reg931_done;
  wire par_done_reg932_in;
  wire par_done_reg932_write_en;
  wire par_done_reg932_clk;
  wire par_done_reg932_out;
  wire par_done_reg932_done;
  wire par_done_reg933_in;
  wire par_done_reg933_write_en;
  wire par_done_reg933_clk;
  wire par_done_reg933_out;
  wire par_done_reg933_done;
  wire par_done_reg934_in;
  wire par_done_reg934_write_en;
  wire par_done_reg934_clk;
  wire par_done_reg934_out;
  wire par_done_reg934_done;
  wire par_done_reg935_in;
  wire par_done_reg935_write_en;
  wire par_done_reg935_clk;
  wire par_done_reg935_out;
  wire par_done_reg935_done;
  wire par_done_reg936_in;
  wire par_done_reg936_write_en;
  wire par_done_reg936_clk;
  wire par_done_reg936_out;
  wire par_done_reg936_done;
  wire par_done_reg937_in;
  wire par_done_reg937_write_en;
  wire par_done_reg937_clk;
  wire par_done_reg937_out;
  wire par_done_reg937_done;
  wire par_done_reg938_in;
  wire par_done_reg938_write_en;
  wire par_done_reg938_clk;
  wire par_done_reg938_out;
  wire par_done_reg938_done;
  wire par_done_reg939_in;
  wire par_done_reg939_write_en;
  wire par_done_reg939_clk;
  wire par_done_reg939_out;
  wire par_done_reg939_done;
  wire par_done_reg940_in;
  wire par_done_reg940_write_en;
  wire par_done_reg940_clk;
  wire par_done_reg940_out;
  wire par_done_reg940_done;
  wire par_done_reg941_in;
  wire par_done_reg941_write_en;
  wire par_done_reg941_clk;
  wire par_done_reg941_out;
  wire par_done_reg941_done;
  wire par_done_reg942_in;
  wire par_done_reg942_write_en;
  wire par_done_reg942_clk;
  wire par_done_reg942_out;
  wire par_done_reg942_done;
  wire par_done_reg943_in;
  wire par_done_reg943_write_en;
  wire par_done_reg943_clk;
  wire par_done_reg943_out;
  wire par_done_reg943_done;
  wire par_done_reg944_in;
  wire par_done_reg944_write_en;
  wire par_done_reg944_clk;
  wire par_done_reg944_out;
  wire par_done_reg944_done;
  wire par_done_reg945_in;
  wire par_done_reg945_write_en;
  wire par_done_reg945_clk;
  wire par_done_reg945_out;
  wire par_done_reg945_done;
  wire par_done_reg946_in;
  wire par_done_reg946_write_en;
  wire par_done_reg946_clk;
  wire par_done_reg946_out;
  wire par_done_reg946_done;
  wire par_done_reg947_in;
  wire par_done_reg947_write_en;
  wire par_done_reg947_clk;
  wire par_done_reg947_out;
  wire par_done_reg947_done;
  wire par_done_reg948_in;
  wire par_done_reg948_write_en;
  wire par_done_reg948_clk;
  wire par_done_reg948_out;
  wire par_done_reg948_done;
  wire par_done_reg949_in;
  wire par_done_reg949_write_en;
  wire par_done_reg949_clk;
  wire par_done_reg949_out;
  wire par_done_reg949_done;
  wire par_done_reg950_in;
  wire par_done_reg950_write_en;
  wire par_done_reg950_clk;
  wire par_done_reg950_out;
  wire par_done_reg950_done;
  wire par_done_reg951_in;
  wire par_done_reg951_write_en;
  wire par_done_reg951_clk;
  wire par_done_reg951_out;
  wire par_done_reg951_done;
  wire par_done_reg952_in;
  wire par_done_reg952_write_en;
  wire par_done_reg952_clk;
  wire par_done_reg952_out;
  wire par_done_reg952_done;
  wire par_done_reg953_in;
  wire par_done_reg953_write_en;
  wire par_done_reg953_clk;
  wire par_done_reg953_out;
  wire par_done_reg953_done;
  wire par_done_reg954_in;
  wire par_done_reg954_write_en;
  wire par_done_reg954_clk;
  wire par_done_reg954_out;
  wire par_done_reg954_done;
  wire par_done_reg955_in;
  wire par_done_reg955_write_en;
  wire par_done_reg955_clk;
  wire par_done_reg955_out;
  wire par_done_reg955_done;
  wire par_done_reg956_in;
  wire par_done_reg956_write_en;
  wire par_done_reg956_clk;
  wire par_done_reg956_out;
  wire par_done_reg956_done;
  wire par_done_reg957_in;
  wire par_done_reg957_write_en;
  wire par_done_reg957_clk;
  wire par_done_reg957_out;
  wire par_done_reg957_done;
  wire par_done_reg958_in;
  wire par_done_reg958_write_en;
  wire par_done_reg958_clk;
  wire par_done_reg958_out;
  wire par_done_reg958_done;
  wire par_done_reg959_in;
  wire par_done_reg959_write_en;
  wire par_done_reg959_clk;
  wire par_done_reg959_out;
  wire par_done_reg959_done;
  wire par_done_reg960_in;
  wire par_done_reg960_write_en;
  wire par_done_reg960_clk;
  wire par_done_reg960_out;
  wire par_done_reg960_done;
  wire par_done_reg961_in;
  wire par_done_reg961_write_en;
  wire par_done_reg961_clk;
  wire par_done_reg961_out;
  wire par_done_reg961_done;
  wire par_done_reg962_in;
  wire par_done_reg962_write_en;
  wire par_done_reg962_clk;
  wire par_done_reg962_out;
  wire par_done_reg962_done;
  wire par_done_reg963_in;
  wire par_done_reg963_write_en;
  wire par_done_reg963_clk;
  wire par_done_reg963_out;
  wire par_done_reg963_done;
  wire par_done_reg964_in;
  wire par_done_reg964_write_en;
  wire par_done_reg964_clk;
  wire par_done_reg964_out;
  wire par_done_reg964_done;
  wire par_done_reg965_in;
  wire par_done_reg965_write_en;
  wire par_done_reg965_clk;
  wire par_done_reg965_out;
  wire par_done_reg965_done;
  wire par_done_reg966_in;
  wire par_done_reg966_write_en;
  wire par_done_reg966_clk;
  wire par_done_reg966_out;
  wire par_done_reg966_done;
  wire par_done_reg967_in;
  wire par_done_reg967_write_en;
  wire par_done_reg967_clk;
  wire par_done_reg967_out;
  wire par_done_reg967_done;
  wire par_done_reg968_in;
  wire par_done_reg968_write_en;
  wire par_done_reg968_clk;
  wire par_done_reg968_out;
  wire par_done_reg968_done;
  wire par_done_reg969_in;
  wire par_done_reg969_write_en;
  wire par_done_reg969_clk;
  wire par_done_reg969_out;
  wire par_done_reg969_done;
  wire par_done_reg970_in;
  wire par_done_reg970_write_en;
  wire par_done_reg970_clk;
  wire par_done_reg970_out;
  wire par_done_reg970_done;
  wire par_done_reg971_in;
  wire par_done_reg971_write_en;
  wire par_done_reg971_clk;
  wire par_done_reg971_out;
  wire par_done_reg971_done;
  wire par_done_reg972_in;
  wire par_done_reg972_write_en;
  wire par_done_reg972_clk;
  wire par_done_reg972_out;
  wire par_done_reg972_done;
  wire par_done_reg973_in;
  wire par_done_reg973_write_en;
  wire par_done_reg973_clk;
  wire par_done_reg973_out;
  wire par_done_reg973_done;
  wire par_done_reg974_in;
  wire par_done_reg974_write_en;
  wire par_done_reg974_clk;
  wire par_done_reg974_out;
  wire par_done_reg974_done;
  wire par_done_reg975_in;
  wire par_done_reg975_write_en;
  wire par_done_reg975_clk;
  wire par_done_reg975_out;
  wire par_done_reg975_done;
  wire par_done_reg976_in;
  wire par_done_reg976_write_en;
  wire par_done_reg976_clk;
  wire par_done_reg976_out;
  wire par_done_reg976_done;
  wire par_done_reg977_in;
  wire par_done_reg977_write_en;
  wire par_done_reg977_clk;
  wire par_done_reg977_out;
  wire par_done_reg977_done;
  wire par_done_reg978_in;
  wire par_done_reg978_write_en;
  wire par_done_reg978_clk;
  wire par_done_reg978_out;
  wire par_done_reg978_done;
  wire par_done_reg979_in;
  wire par_done_reg979_write_en;
  wire par_done_reg979_clk;
  wire par_done_reg979_out;
  wire par_done_reg979_done;
  wire par_done_reg980_in;
  wire par_done_reg980_write_en;
  wire par_done_reg980_clk;
  wire par_done_reg980_out;
  wire par_done_reg980_done;
  wire par_done_reg981_in;
  wire par_done_reg981_write_en;
  wire par_done_reg981_clk;
  wire par_done_reg981_out;
  wire par_done_reg981_done;
  wire par_done_reg982_in;
  wire par_done_reg982_write_en;
  wire par_done_reg982_clk;
  wire par_done_reg982_out;
  wire par_done_reg982_done;
  wire par_done_reg983_in;
  wire par_done_reg983_write_en;
  wire par_done_reg983_clk;
  wire par_done_reg983_out;
  wire par_done_reg983_done;
  wire par_done_reg984_in;
  wire par_done_reg984_write_en;
  wire par_done_reg984_clk;
  wire par_done_reg984_out;
  wire par_done_reg984_done;
  wire par_done_reg985_in;
  wire par_done_reg985_write_en;
  wire par_done_reg985_clk;
  wire par_done_reg985_out;
  wire par_done_reg985_done;
  wire par_done_reg986_in;
  wire par_done_reg986_write_en;
  wire par_done_reg986_clk;
  wire par_done_reg986_out;
  wire par_done_reg986_done;
  wire par_done_reg987_in;
  wire par_done_reg987_write_en;
  wire par_done_reg987_clk;
  wire par_done_reg987_out;
  wire par_done_reg987_done;
  wire par_done_reg988_in;
  wire par_done_reg988_write_en;
  wire par_done_reg988_clk;
  wire par_done_reg988_out;
  wire par_done_reg988_done;
  wire par_done_reg989_in;
  wire par_done_reg989_write_en;
  wire par_done_reg989_clk;
  wire par_done_reg989_out;
  wire par_done_reg989_done;
  wire par_done_reg990_in;
  wire par_done_reg990_write_en;
  wire par_done_reg990_clk;
  wire par_done_reg990_out;
  wire par_done_reg990_done;
  wire par_done_reg991_in;
  wire par_done_reg991_write_en;
  wire par_done_reg991_clk;
  wire par_done_reg991_out;
  wire par_done_reg991_done;
  wire par_done_reg992_in;
  wire par_done_reg992_write_en;
  wire par_done_reg992_clk;
  wire par_done_reg992_out;
  wire par_done_reg992_done;
  wire par_done_reg993_in;
  wire par_done_reg993_write_en;
  wire par_done_reg993_clk;
  wire par_done_reg993_out;
  wire par_done_reg993_done;
  wire par_done_reg994_in;
  wire par_done_reg994_write_en;
  wire par_done_reg994_clk;
  wire par_done_reg994_out;
  wire par_done_reg994_done;
  wire par_done_reg995_in;
  wire par_done_reg995_write_en;
  wire par_done_reg995_clk;
  wire par_done_reg995_out;
  wire par_done_reg995_done;
  wire par_reset25_in;
  wire par_reset25_write_en;
  wire par_reset25_clk;
  wire par_reset25_out;
  wire par_reset25_done;
  wire par_done_reg996_in;
  wire par_done_reg996_write_en;
  wire par_done_reg996_clk;
  wire par_done_reg996_out;
  wire par_done_reg996_done;
  wire par_done_reg997_in;
  wire par_done_reg997_write_en;
  wire par_done_reg997_clk;
  wire par_done_reg997_out;
  wire par_done_reg997_done;
  wire par_done_reg998_in;
  wire par_done_reg998_write_en;
  wire par_done_reg998_clk;
  wire par_done_reg998_out;
  wire par_done_reg998_done;
  wire par_done_reg999_in;
  wire par_done_reg999_write_en;
  wire par_done_reg999_clk;
  wire par_done_reg999_out;
  wire par_done_reg999_done;
  wire par_done_reg1000_in;
  wire par_done_reg1000_write_en;
  wire par_done_reg1000_clk;
  wire par_done_reg1000_out;
  wire par_done_reg1000_done;
  wire par_done_reg1001_in;
  wire par_done_reg1001_write_en;
  wire par_done_reg1001_clk;
  wire par_done_reg1001_out;
  wire par_done_reg1001_done;
  wire par_done_reg1002_in;
  wire par_done_reg1002_write_en;
  wire par_done_reg1002_clk;
  wire par_done_reg1002_out;
  wire par_done_reg1002_done;
  wire par_done_reg1003_in;
  wire par_done_reg1003_write_en;
  wire par_done_reg1003_clk;
  wire par_done_reg1003_out;
  wire par_done_reg1003_done;
  wire par_done_reg1004_in;
  wire par_done_reg1004_write_en;
  wire par_done_reg1004_clk;
  wire par_done_reg1004_out;
  wire par_done_reg1004_done;
  wire par_done_reg1005_in;
  wire par_done_reg1005_write_en;
  wire par_done_reg1005_clk;
  wire par_done_reg1005_out;
  wire par_done_reg1005_done;
  wire par_done_reg1006_in;
  wire par_done_reg1006_write_en;
  wire par_done_reg1006_clk;
  wire par_done_reg1006_out;
  wire par_done_reg1006_done;
  wire par_done_reg1007_in;
  wire par_done_reg1007_write_en;
  wire par_done_reg1007_clk;
  wire par_done_reg1007_out;
  wire par_done_reg1007_done;
  wire par_done_reg1008_in;
  wire par_done_reg1008_write_en;
  wire par_done_reg1008_clk;
  wire par_done_reg1008_out;
  wire par_done_reg1008_done;
  wire par_done_reg1009_in;
  wire par_done_reg1009_write_en;
  wire par_done_reg1009_clk;
  wire par_done_reg1009_out;
  wire par_done_reg1009_done;
  wire par_done_reg1010_in;
  wire par_done_reg1010_write_en;
  wire par_done_reg1010_clk;
  wire par_done_reg1010_out;
  wire par_done_reg1010_done;
  wire par_done_reg1011_in;
  wire par_done_reg1011_write_en;
  wire par_done_reg1011_clk;
  wire par_done_reg1011_out;
  wire par_done_reg1011_done;
  wire par_done_reg1012_in;
  wire par_done_reg1012_write_en;
  wire par_done_reg1012_clk;
  wire par_done_reg1012_out;
  wire par_done_reg1012_done;
  wire par_done_reg1013_in;
  wire par_done_reg1013_write_en;
  wire par_done_reg1013_clk;
  wire par_done_reg1013_out;
  wire par_done_reg1013_done;
  wire par_done_reg1014_in;
  wire par_done_reg1014_write_en;
  wire par_done_reg1014_clk;
  wire par_done_reg1014_out;
  wire par_done_reg1014_done;
  wire par_done_reg1015_in;
  wire par_done_reg1015_write_en;
  wire par_done_reg1015_clk;
  wire par_done_reg1015_out;
  wire par_done_reg1015_done;
  wire par_done_reg1016_in;
  wire par_done_reg1016_write_en;
  wire par_done_reg1016_clk;
  wire par_done_reg1016_out;
  wire par_done_reg1016_done;
  wire par_done_reg1017_in;
  wire par_done_reg1017_write_en;
  wire par_done_reg1017_clk;
  wire par_done_reg1017_out;
  wire par_done_reg1017_done;
  wire par_done_reg1018_in;
  wire par_done_reg1018_write_en;
  wire par_done_reg1018_clk;
  wire par_done_reg1018_out;
  wire par_done_reg1018_done;
  wire par_done_reg1019_in;
  wire par_done_reg1019_write_en;
  wire par_done_reg1019_clk;
  wire par_done_reg1019_out;
  wire par_done_reg1019_done;
  wire par_done_reg1020_in;
  wire par_done_reg1020_write_en;
  wire par_done_reg1020_clk;
  wire par_done_reg1020_out;
  wire par_done_reg1020_done;
  wire par_done_reg1021_in;
  wire par_done_reg1021_write_en;
  wire par_done_reg1021_clk;
  wire par_done_reg1021_out;
  wire par_done_reg1021_done;
  wire par_done_reg1022_in;
  wire par_done_reg1022_write_en;
  wire par_done_reg1022_clk;
  wire par_done_reg1022_out;
  wire par_done_reg1022_done;
  wire par_done_reg1023_in;
  wire par_done_reg1023_write_en;
  wire par_done_reg1023_clk;
  wire par_done_reg1023_out;
  wire par_done_reg1023_done;
  wire par_done_reg1024_in;
  wire par_done_reg1024_write_en;
  wire par_done_reg1024_clk;
  wire par_done_reg1024_out;
  wire par_done_reg1024_done;
  wire par_done_reg1025_in;
  wire par_done_reg1025_write_en;
  wire par_done_reg1025_clk;
  wire par_done_reg1025_out;
  wire par_done_reg1025_done;
  wire par_done_reg1026_in;
  wire par_done_reg1026_write_en;
  wire par_done_reg1026_clk;
  wire par_done_reg1026_out;
  wire par_done_reg1026_done;
  wire par_done_reg1027_in;
  wire par_done_reg1027_write_en;
  wire par_done_reg1027_clk;
  wire par_done_reg1027_out;
  wire par_done_reg1027_done;
  wire par_done_reg1028_in;
  wire par_done_reg1028_write_en;
  wire par_done_reg1028_clk;
  wire par_done_reg1028_out;
  wire par_done_reg1028_done;
  wire par_done_reg1029_in;
  wire par_done_reg1029_write_en;
  wire par_done_reg1029_clk;
  wire par_done_reg1029_out;
  wire par_done_reg1029_done;
  wire par_done_reg1030_in;
  wire par_done_reg1030_write_en;
  wire par_done_reg1030_clk;
  wire par_done_reg1030_out;
  wire par_done_reg1030_done;
  wire par_done_reg1031_in;
  wire par_done_reg1031_write_en;
  wire par_done_reg1031_clk;
  wire par_done_reg1031_out;
  wire par_done_reg1031_done;
  wire par_done_reg1032_in;
  wire par_done_reg1032_write_en;
  wire par_done_reg1032_clk;
  wire par_done_reg1032_out;
  wire par_done_reg1032_done;
  wire par_done_reg1033_in;
  wire par_done_reg1033_write_en;
  wire par_done_reg1033_clk;
  wire par_done_reg1033_out;
  wire par_done_reg1033_done;
  wire par_done_reg1034_in;
  wire par_done_reg1034_write_en;
  wire par_done_reg1034_clk;
  wire par_done_reg1034_out;
  wire par_done_reg1034_done;
  wire par_done_reg1035_in;
  wire par_done_reg1035_write_en;
  wire par_done_reg1035_clk;
  wire par_done_reg1035_out;
  wire par_done_reg1035_done;
  wire par_done_reg1036_in;
  wire par_done_reg1036_write_en;
  wire par_done_reg1036_clk;
  wire par_done_reg1036_out;
  wire par_done_reg1036_done;
  wire par_done_reg1037_in;
  wire par_done_reg1037_write_en;
  wire par_done_reg1037_clk;
  wire par_done_reg1037_out;
  wire par_done_reg1037_done;
  wire par_done_reg1038_in;
  wire par_done_reg1038_write_en;
  wire par_done_reg1038_clk;
  wire par_done_reg1038_out;
  wire par_done_reg1038_done;
  wire par_done_reg1039_in;
  wire par_done_reg1039_write_en;
  wire par_done_reg1039_clk;
  wire par_done_reg1039_out;
  wire par_done_reg1039_done;
  wire par_done_reg1040_in;
  wire par_done_reg1040_write_en;
  wire par_done_reg1040_clk;
  wire par_done_reg1040_out;
  wire par_done_reg1040_done;
  wire par_done_reg1041_in;
  wire par_done_reg1041_write_en;
  wire par_done_reg1041_clk;
  wire par_done_reg1041_out;
  wire par_done_reg1041_done;
  wire par_done_reg1042_in;
  wire par_done_reg1042_write_en;
  wire par_done_reg1042_clk;
  wire par_done_reg1042_out;
  wire par_done_reg1042_done;
  wire par_done_reg1043_in;
  wire par_done_reg1043_write_en;
  wire par_done_reg1043_clk;
  wire par_done_reg1043_out;
  wire par_done_reg1043_done;
  wire par_done_reg1044_in;
  wire par_done_reg1044_write_en;
  wire par_done_reg1044_clk;
  wire par_done_reg1044_out;
  wire par_done_reg1044_done;
  wire par_done_reg1045_in;
  wire par_done_reg1045_write_en;
  wire par_done_reg1045_clk;
  wire par_done_reg1045_out;
  wire par_done_reg1045_done;
  wire par_done_reg1046_in;
  wire par_done_reg1046_write_en;
  wire par_done_reg1046_clk;
  wire par_done_reg1046_out;
  wire par_done_reg1046_done;
  wire par_done_reg1047_in;
  wire par_done_reg1047_write_en;
  wire par_done_reg1047_clk;
  wire par_done_reg1047_out;
  wire par_done_reg1047_done;
  wire par_done_reg1048_in;
  wire par_done_reg1048_write_en;
  wire par_done_reg1048_clk;
  wire par_done_reg1048_out;
  wire par_done_reg1048_done;
  wire par_done_reg1049_in;
  wire par_done_reg1049_write_en;
  wire par_done_reg1049_clk;
  wire par_done_reg1049_out;
  wire par_done_reg1049_done;
  wire par_reset26_in;
  wire par_reset26_write_en;
  wire par_reset26_clk;
  wire par_reset26_out;
  wire par_reset26_done;
  wire par_done_reg1050_in;
  wire par_done_reg1050_write_en;
  wire par_done_reg1050_clk;
  wire par_done_reg1050_out;
  wire par_done_reg1050_done;
  wire par_done_reg1051_in;
  wire par_done_reg1051_write_en;
  wire par_done_reg1051_clk;
  wire par_done_reg1051_out;
  wire par_done_reg1051_done;
  wire par_done_reg1052_in;
  wire par_done_reg1052_write_en;
  wire par_done_reg1052_clk;
  wire par_done_reg1052_out;
  wire par_done_reg1052_done;
  wire par_done_reg1053_in;
  wire par_done_reg1053_write_en;
  wire par_done_reg1053_clk;
  wire par_done_reg1053_out;
  wire par_done_reg1053_done;
  wire par_done_reg1054_in;
  wire par_done_reg1054_write_en;
  wire par_done_reg1054_clk;
  wire par_done_reg1054_out;
  wire par_done_reg1054_done;
  wire par_done_reg1055_in;
  wire par_done_reg1055_write_en;
  wire par_done_reg1055_clk;
  wire par_done_reg1055_out;
  wire par_done_reg1055_done;
  wire par_done_reg1056_in;
  wire par_done_reg1056_write_en;
  wire par_done_reg1056_clk;
  wire par_done_reg1056_out;
  wire par_done_reg1056_done;
  wire par_done_reg1057_in;
  wire par_done_reg1057_write_en;
  wire par_done_reg1057_clk;
  wire par_done_reg1057_out;
  wire par_done_reg1057_done;
  wire par_done_reg1058_in;
  wire par_done_reg1058_write_en;
  wire par_done_reg1058_clk;
  wire par_done_reg1058_out;
  wire par_done_reg1058_done;
  wire par_done_reg1059_in;
  wire par_done_reg1059_write_en;
  wire par_done_reg1059_clk;
  wire par_done_reg1059_out;
  wire par_done_reg1059_done;
  wire par_done_reg1060_in;
  wire par_done_reg1060_write_en;
  wire par_done_reg1060_clk;
  wire par_done_reg1060_out;
  wire par_done_reg1060_done;
  wire par_done_reg1061_in;
  wire par_done_reg1061_write_en;
  wire par_done_reg1061_clk;
  wire par_done_reg1061_out;
  wire par_done_reg1061_done;
  wire par_done_reg1062_in;
  wire par_done_reg1062_write_en;
  wire par_done_reg1062_clk;
  wire par_done_reg1062_out;
  wire par_done_reg1062_done;
  wire par_done_reg1063_in;
  wire par_done_reg1063_write_en;
  wire par_done_reg1063_clk;
  wire par_done_reg1063_out;
  wire par_done_reg1063_done;
  wire par_done_reg1064_in;
  wire par_done_reg1064_write_en;
  wire par_done_reg1064_clk;
  wire par_done_reg1064_out;
  wire par_done_reg1064_done;
  wire par_done_reg1065_in;
  wire par_done_reg1065_write_en;
  wire par_done_reg1065_clk;
  wire par_done_reg1065_out;
  wire par_done_reg1065_done;
  wire par_done_reg1066_in;
  wire par_done_reg1066_write_en;
  wire par_done_reg1066_clk;
  wire par_done_reg1066_out;
  wire par_done_reg1066_done;
  wire par_done_reg1067_in;
  wire par_done_reg1067_write_en;
  wire par_done_reg1067_clk;
  wire par_done_reg1067_out;
  wire par_done_reg1067_done;
  wire par_done_reg1068_in;
  wire par_done_reg1068_write_en;
  wire par_done_reg1068_clk;
  wire par_done_reg1068_out;
  wire par_done_reg1068_done;
  wire par_done_reg1069_in;
  wire par_done_reg1069_write_en;
  wire par_done_reg1069_clk;
  wire par_done_reg1069_out;
  wire par_done_reg1069_done;
  wire par_done_reg1070_in;
  wire par_done_reg1070_write_en;
  wire par_done_reg1070_clk;
  wire par_done_reg1070_out;
  wire par_done_reg1070_done;
  wire par_done_reg1071_in;
  wire par_done_reg1071_write_en;
  wire par_done_reg1071_clk;
  wire par_done_reg1071_out;
  wire par_done_reg1071_done;
  wire par_done_reg1072_in;
  wire par_done_reg1072_write_en;
  wire par_done_reg1072_clk;
  wire par_done_reg1072_out;
  wire par_done_reg1072_done;
  wire par_done_reg1073_in;
  wire par_done_reg1073_write_en;
  wire par_done_reg1073_clk;
  wire par_done_reg1073_out;
  wire par_done_reg1073_done;
  wire par_done_reg1074_in;
  wire par_done_reg1074_write_en;
  wire par_done_reg1074_clk;
  wire par_done_reg1074_out;
  wire par_done_reg1074_done;
  wire par_done_reg1075_in;
  wire par_done_reg1075_write_en;
  wire par_done_reg1075_clk;
  wire par_done_reg1075_out;
  wire par_done_reg1075_done;
  wire par_done_reg1076_in;
  wire par_done_reg1076_write_en;
  wire par_done_reg1076_clk;
  wire par_done_reg1076_out;
  wire par_done_reg1076_done;
  wire par_done_reg1077_in;
  wire par_done_reg1077_write_en;
  wire par_done_reg1077_clk;
  wire par_done_reg1077_out;
  wire par_done_reg1077_done;
  wire par_done_reg1078_in;
  wire par_done_reg1078_write_en;
  wire par_done_reg1078_clk;
  wire par_done_reg1078_out;
  wire par_done_reg1078_done;
  wire par_done_reg1079_in;
  wire par_done_reg1079_write_en;
  wire par_done_reg1079_clk;
  wire par_done_reg1079_out;
  wire par_done_reg1079_done;
  wire par_done_reg1080_in;
  wire par_done_reg1080_write_en;
  wire par_done_reg1080_clk;
  wire par_done_reg1080_out;
  wire par_done_reg1080_done;
  wire par_done_reg1081_in;
  wire par_done_reg1081_write_en;
  wire par_done_reg1081_clk;
  wire par_done_reg1081_out;
  wire par_done_reg1081_done;
  wire par_done_reg1082_in;
  wire par_done_reg1082_write_en;
  wire par_done_reg1082_clk;
  wire par_done_reg1082_out;
  wire par_done_reg1082_done;
  wire par_done_reg1083_in;
  wire par_done_reg1083_write_en;
  wire par_done_reg1083_clk;
  wire par_done_reg1083_out;
  wire par_done_reg1083_done;
  wire par_done_reg1084_in;
  wire par_done_reg1084_write_en;
  wire par_done_reg1084_clk;
  wire par_done_reg1084_out;
  wire par_done_reg1084_done;
  wire par_done_reg1085_in;
  wire par_done_reg1085_write_en;
  wire par_done_reg1085_clk;
  wire par_done_reg1085_out;
  wire par_done_reg1085_done;
  wire par_done_reg1086_in;
  wire par_done_reg1086_write_en;
  wire par_done_reg1086_clk;
  wire par_done_reg1086_out;
  wire par_done_reg1086_done;
  wire par_done_reg1087_in;
  wire par_done_reg1087_write_en;
  wire par_done_reg1087_clk;
  wire par_done_reg1087_out;
  wire par_done_reg1087_done;
  wire par_done_reg1088_in;
  wire par_done_reg1088_write_en;
  wire par_done_reg1088_clk;
  wire par_done_reg1088_out;
  wire par_done_reg1088_done;
  wire par_done_reg1089_in;
  wire par_done_reg1089_write_en;
  wire par_done_reg1089_clk;
  wire par_done_reg1089_out;
  wire par_done_reg1089_done;
  wire par_done_reg1090_in;
  wire par_done_reg1090_write_en;
  wire par_done_reg1090_clk;
  wire par_done_reg1090_out;
  wire par_done_reg1090_done;
  wire par_done_reg1091_in;
  wire par_done_reg1091_write_en;
  wire par_done_reg1091_clk;
  wire par_done_reg1091_out;
  wire par_done_reg1091_done;
  wire par_done_reg1092_in;
  wire par_done_reg1092_write_en;
  wire par_done_reg1092_clk;
  wire par_done_reg1092_out;
  wire par_done_reg1092_done;
  wire par_done_reg1093_in;
  wire par_done_reg1093_write_en;
  wire par_done_reg1093_clk;
  wire par_done_reg1093_out;
  wire par_done_reg1093_done;
  wire par_done_reg1094_in;
  wire par_done_reg1094_write_en;
  wire par_done_reg1094_clk;
  wire par_done_reg1094_out;
  wire par_done_reg1094_done;
  wire par_done_reg1095_in;
  wire par_done_reg1095_write_en;
  wire par_done_reg1095_clk;
  wire par_done_reg1095_out;
  wire par_done_reg1095_done;
  wire par_done_reg1096_in;
  wire par_done_reg1096_write_en;
  wire par_done_reg1096_clk;
  wire par_done_reg1096_out;
  wire par_done_reg1096_done;
  wire par_done_reg1097_in;
  wire par_done_reg1097_write_en;
  wire par_done_reg1097_clk;
  wire par_done_reg1097_out;
  wire par_done_reg1097_done;
  wire par_done_reg1098_in;
  wire par_done_reg1098_write_en;
  wire par_done_reg1098_clk;
  wire par_done_reg1098_out;
  wire par_done_reg1098_done;
  wire par_done_reg1099_in;
  wire par_done_reg1099_write_en;
  wire par_done_reg1099_clk;
  wire par_done_reg1099_out;
  wire par_done_reg1099_done;
  wire par_done_reg1100_in;
  wire par_done_reg1100_write_en;
  wire par_done_reg1100_clk;
  wire par_done_reg1100_out;
  wire par_done_reg1100_done;
  wire par_done_reg1101_in;
  wire par_done_reg1101_write_en;
  wire par_done_reg1101_clk;
  wire par_done_reg1101_out;
  wire par_done_reg1101_done;
  wire par_done_reg1102_in;
  wire par_done_reg1102_write_en;
  wire par_done_reg1102_clk;
  wire par_done_reg1102_out;
  wire par_done_reg1102_done;
  wire par_done_reg1103_in;
  wire par_done_reg1103_write_en;
  wire par_done_reg1103_clk;
  wire par_done_reg1103_out;
  wire par_done_reg1103_done;
  wire par_done_reg1104_in;
  wire par_done_reg1104_write_en;
  wire par_done_reg1104_clk;
  wire par_done_reg1104_out;
  wire par_done_reg1104_done;
  wire par_done_reg1105_in;
  wire par_done_reg1105_write_en;
  wire par_done_reg1105_clk;
  wire par_done_reg1105_out;
  wire par_done_reg1105_done;
  wire par_done_reg1106_in;
  wire par_done_reg1106_write_en;
  wire par_done_reg1106_clk;
  wire par_done_reg1106_out;
  wire par_done_reg1106_done;
  wire par_done_reg1107_in;
  wire par_done_reg1107_write_en;
  wire par_done_reg1107_clk;
  wire par_done_reg1107_out;
  wire par_done_reg1107_done;
  wire par_done_reg1108_in;
  wire par_done_reg1108_write_en;
  wire par_done_reg1108_clk;
  wire par_done_reg1108_out;
  wire par_done_reg1108_done;
  wire par_done_reg1109_in;
  wire par_done_reg1109_write_en;
  wire par_done_reg1109_clk;
  wire par_done_reg1109_out;
  wire par_done_reg1109_done;
  wire par_done_reg1110_in;
  wire par_done_reg1110_write_en;
  wire par_done_reg1110_clk;
  wire par_done_reg1110_out;
  wire par_done_reg1110_done;
  wire par_done_reg1111_in;
  wire par_done_reg1111_write_en;
  wire par_done_reg1111_clk;
  wire par_done_reg1111_out;
  wire par_done_reg1111_done;
  wire par_done_reg1112_in;
  wire par_done_reg1112_write_en;
  wire par_done_reg1112_clk;
  wire par_done_reg1112_out;
  wire par_done_reg1112_done;
  wire par_done_reg1113_in;
  wire par_done_reg1113_write_en;
  wire par_done_reg1113_clk;
  wire par_done_reg1113_out;
  wire par_done_reg1113_done;
  wire par_done_reg1114_in;
  wire par_done_reg1114_write_en;
  wire par_done_reg1114_clk;
  wire par_done_reg1114_out;
  wire par_done_reg1114_done;
  wire par_done_reg1115_in;
  wire par_done_reg1115_write_en;
  wire par_done_reg1115_clk;
  wire par_done_reg1115_out;
  wire par_done_reg1115_done;
  wire par_done_reg1116_in;
  wire par_done_reg1116_write_en;
  wire par_done_reg1116_clk;
  wire par_done_reg1116_out;
  wire par_done_reg1116_done;
  wire par_done_reg1117_in;
  wire par_done_reg1117_write_en;
  wire par_done_reg1117_clk;
  wire par_done_reg1117_out;
  wire par_done_reg1117_done;
  wire par_done_reg1118_in;
  wire par_done_reg1118_write_en;
  wire par_done_reg1118_clk;
  wire par_done_reg1118_out;
  wire par_done_reg1118_done;
  wire par_done_reg1119_in;
  wire par_done_reg1119_write_en;
  wire par_done_reg1119_clk;
  wire par_done_reg1119_out;
  wire par_done_reg1119_done;
  wire par_done_reg1120_in;
  wire par_done_reg1120_write_en;
  wire par_done_reg1120_clk;
  wire par_done_reg1120_out;
  wire par_done_reg1120_done;
  wire par_done_reg1121_in;
  wire par_done_reg1121_write_en;
  wire par_done_reg1121_clk;
  wire par_done_reg1121_out;
  wire par_done_reg1121_done;
  wire par_done_reg1122_in;
  wire par_done_reg1122_write_en;
  wire par_done_reg1122_clk;
  wire par_done_reg1122_out;
  wire par_done_reg1122_done;
  wire par_done_reg1123_in;
  wire par_done_reg1123_write_en;
  wire par_done_reg1123_clk;
  wire par_done_reg1123_out;
  wire par_done_reg1123_done;
  wire par_done_reg1124_in;
  wire par_done_reg1124_write_en;
  wire par_done_reg1124_clk;
  wire par_done_reg1124_out;
  wire par_done_reg1124_done;
  wire par_done_reg1125_in;
  wire par_done_reg1125_write_en;
  wire par_done_reg1125_clk;
  wire par_done_reg1125_out;
  wire par_done_reg1125_done;
  wire par_done_reg1126_in;
  wire par_done_reg1126_write_en;
  wire par_done_reg1126_clk;
  wire par_done_reg1126_out;
  wire par_done_reg1126_done;
  wire par_done_reg1127_in;
  wire par_done_reg1127_write_en;
  wire par_done_reg1127_clk;
  wire par_done_reg1127_out;
  wire par_done_reg1127_done;
  wire par_done_reg1128_in;
  wire par_done_reg1128_write_en;
  wire par_done_reg1128_clk;
  wire par_done_reg1128_out;
  wire par_done_reg1128_done;
  wire par_done_reg1129_in;
  wire par_done_reg1129_write_en;
  wire par_done_reg1129_clk;
  wire par_done_reg1129_out;
  wire par_done_reg1129_done;
  wire par_done_reg1130_in;
  wire par_done_reg1130_write_en;
  wire par_done_reg1130_clk;
  wire par_done_reg1130_out;
  wire par_done_reg1130_done;
  wire par_done_reg1131_in;
  wire par_done_reg1131_write_en;
  wire par_done_reg1131_clk;
  wire par_done_reg1131_out;
  wire par_done_reg1131_done;
  wire par_done_reg1132_in;
  wire par_done_reg1132_write_en;
  wire par_done_reg1132_clk;
  wire par_done_reg1132_out;
  wire par_done_reg1132_done;
  wire par_done_reg1133_in;
  wire par_done_reg1133_write_en;
  wire par_done_reg1133_clk;
  wire par_done_reg1133_out;
  wire par_done_reg1133_done;
  wire par_done_reg1134_in;
  wire par_done_reg1134_write_en;
  wire par_done_reg1134_clk;
  wire par_done_reg1134_out;
  wire par_done_reg1134_done;
  wire par_done_reg1135_in;
  wire par_done_reg1135_write_en;
  wire par_done_reg1135_clk;
  wire par_done_reg1135_out;
  wire par_done_reg1135_done;
  wire par_done_reg1136_in;
  wire par_done_reg1136_write_en;
  wire par_done_reg1136_clk;
  wire par_done_reg1136_out;
  wire par_done_reg1136_done;
  wire par_done_reg1137_in;
  wire par_done_reg1137_write_en;
  wire par_done_reg1137_clk;
  wire par_done_reg1137_out;
  wire par_done_reg1137_done;
  wire par_done_reg1138_in;
  wire par_done_reg1138_write_en;
  wire par_done_reg1138_clk;
  wire par_done_reg1138_out;
  wire par_done_reg1138_done;
  wire par_done_reg1139_in;
  wire par_done_reg1139_write_en;
  wire par_done_reg1139_clk;
  wire par_done_reg1139_out;
  wire par_done_reg1139_done;
  wire par_done_reg1140_in;
  wire par_done_reg1140_write_en;
  wire par_done_reg1140_clk;
  wire par_done_reg1140_out;
  wire par_done_reg1140_done;
  wire par_done_reg1141_in;
  wire par_done_reg1141_write_en;
  wire par_done_reg1141_clk;
  wire par_done_reg1141_out;
  wire par_done_reg1141_done;
  wire par_reset27_in;
  wire par_reset27_write_en;
  wire par_reset27_clk;
  wire par_reset27_out;
  wire par_reset27_done;
  wire par_done_reg1142_in;
  wire par_done_reg1142_write_en;
  wire par_done_reg1142_clk;
  wire par_done_reg1142_out;
  wire par_done_reg1142_done;
  wire par_done_reg1143_in;
  wire par_done_reg1143_write_en;
  wire par_done_reg1143_clk;
  wire par_done_reg1143_out;
  wire par_done_reg1143_done;
  wire par_done_reg1144_in;
  wire par_done_reg1144_write_en;
  wire par_done_reg1144_clk;
  wire par_done_reg1144_out;
  wire par_done_reg1144_done;
  wire par_done_reg1145_in;
  wire par_done_reg1145_write_en;
  wire par_done_reg1145_clk;
  wire par_done_reg1145_out;
  wire par_done_reg1145_done;
  wire par_done_reg1146_in;
  wire par_done_reg1146_write_en;
  wire par_done_reg1146_clk;
  wire par_done_reg1146_out;
  wire par_done_reg1146_done;
  wire par_done_reg1147_in;
  wire par_done_reg1147_write_en;
  wire par_done_reg1147_clk;
  wire par_done_reg1147_out;
  wire par_done_reg1147_done;
  wire par_done_reg1148_in;
  wire par_done_reg1148_write_en;
  wire par_done_reg1148_clk;
  wire par_done_reg1148_out;
  wire par_done_reg1148_done;
  wire par_done_reg1149_in;
  wire par_done_reg1149_write_en;
  wire par_done_reg1149_clk;
  wire par_done_reg1149_out;
  wire par_done_reg1149_done;
  wire par_done_reg1150_in;
  wire par_done_reg1150_write_en;
  wire par_done_reg1150_clk;
  wire par_done_reg1150_out;
  wire par_done_reg1150_done;
  wire par_done_reg1151_in;
  wire par_done_reg1151_write_en;
  wire par_done_reg1151_clk;
  wire par_done_reg1151_out;
  wire par_done_reg1151_done;
  wire par_done_reg1152_in;
  wire par_done_reg1152_write_en;
  wire par_done_reg1152_clk;
  wire par_done_reg1152_out;
  wire par_done_reg1152_done;
  wire par_done_reg1153_in;
  wire par_done_reg1153_write_en;
  wire par_done_reg1153_clk;
  wire par_done_reg1153_out;
  wire par_done_reg1153_done;
  wire par_done_reg1154_in;
  wire par_done_reg1154_write_en;
  wire par_done_reg1154_clk;
  wire par_done_reg1154_out;
  wire par_done_reg1154_done;
  wire par_done_reg1155_in;
  wire par_done_reg1155_write_en;
  wire par_done_reg1155_clk;
  wire par_done_reg1155_out;
  wire par_done_reg1155_done;
  wire par_done_reg1156_in;
  wire par_done_reg1156_write_en;
  wire par_done_reg1156_clk;
  wire par_done_reg1156_out;
  wire par_done_reg1156_done;
  wire par_done_reg1157_in;
  wire par_done_reg1157_write_en;
  wire par_done_reg1157_clk;
  wire par_done_reg1157_out;
  wire par_done_reg1157_done;
  wire par_done_reg1158_in;
  wire par_done_reg1158_write_en;
  wire par_done_reg1158_clk;
  wire par_done_reg1158_out;
  wire par_done_reg1158_done;
  wire par_done_reg1159_in;
  wire par_done_reg1159_write_en;
  wire par_done_reg1159_clk;
  wire par_done_reg1159_out;
  wire par_done_reg1159_done;
  wire par_done_reg1160_in;
  wire par_done_reg1160_write_en;
  wire par_done_reg1160_clk;
  wire par_done_reg1160_out;
  wire par_done_reg1160_done;
  wire par_done_reg1161_in;
  wire par_done_reg1161_write_en;
  wire par_done_reg1161_clk;
  wire par_done_reg1161_out;
  wire par_done_reg1161_done;
  wire par_done_reg1162_in;
  wire par_done_reg1162_write_en;
  wire par_done_reg1162_clk;
  wire par_done_reg1162_out;
  wire par_done_reg1162_done;
  wire par_done_reg1163_in;
  wire par_done_reg1163_write_en;
  wire par_done_reg1163_clk;
  wire par_done_reg1163_out;
  wire par_done_reg1163_done;
  wire par_done_reg1164_in;
  wire par_done_reg1164_write_en;
  wire par_done_reg1164_clk;
  wire par_done_reg1164_out;
  wire par_done_reg1164_done;
  wire par_done_reg1165_in;
  wire par_done_reg1165_write_en;
  wire par_done_reg1165_clk;
  wire par_done_reg1165_out;
  wire par_done_reg1165_done;
  wire par_done_reg1166_in;
  wire par_done_reg1166_write_en;
  wire par_done_reg1166_clk;
  wire par_done_reg1166_out;
  wire par_done_reg1166_done;
  wire par_done_reg1167_in;
  wire par_done_reg1167_write_en;
  wire par_done_reg1167_clk;
  wire par_done_reg1167_out;
  wire par_done_reg1167_done;
  wire par_done_reg1168_in;
  wire par_done_reg1168_write_en;
  wire par_done_reg1168_clk;
  wire par_done_reg1168_out;
  wire par_done_reg1168_done;
  wire par_done_reg1169_in;
  wire par_done_reg1169_write_en;
  wire par_done_reg1169_clk;
  wire par_done_reg1169_out;
  wire par_done_reg1169_done;
  wire par_done_reg1170_in;
  wire par_done_reg1170_write_en;
  wire par_done_reg1170_clk;
  wire par_done_reg1170_out;
  wire par_done_reg1170_done;
  wire par_done_reg1171_in;
  wire par_done_reg1171_write_en;
  wire par_done_reg1171_clk;
  wire par_done_reg1171_out;
  wire par_done_reg1171_done;
  wire par_done_reg1172_in;
  wire par_done_reg1172_write_en;
  wire par_done_reg1172_clk;
  wire par_done_reg1172_out;
  wire par_done_reg1172_done;
  wire par_done_reg1173_in;
  wire par_done_reg1173_write_en;
  wire par_done_reg1173_clk;
  wire par_done_reg1173_out;
  wire par_done_reg1173_done;
  wire par_done_reg1174_in;
  wire par_done_reg1174_write_en;
  wire par_done_reg1174_clk;
  wire par_done_reg1174_out;
  wire par_done_reg1174_done;
  wire par_done_reg1175_in;
  wire par_done_reg1175_write_en;
  wire par_done_reg1175_clk;
  wire par_done_reg1175_out;
  wire par_done_reg1175_done;
  wire par_done_reg1176_in;
  wire par_done_reg1176_write_en;
  wire par_done_reg1176_clk;
  wire par_done_reg1176_out;
  wire par_done_reg1176_done;
  wire par_done_reg1177_in;
  wire par_done_reg1177_write_en;
  wire par_done_reg1177_clk;
  wire par_done_reg1177_out;
  wire par_done_reg1177_done;
  wire par_done_reg1178_in;
  wire par_done_reg1178_write_en;
  wire par_done_reg1178_clk;
  wire par_done_reg1178_out;
  wire par_done_reg1178_done;
  wire par_done_reg1179_in;
  wire par_done_reg1179_write_en;
  wire par_done_reg1179_clk;
  wire par_done_reg1179_out;
  wire par_done_reg1179_done;
  wire par_done_reg1180_in;
  wire par_done_reg1180_write_en;
  wire par_done_reg1180_clk;
  wire par_done_reg1180_out;
  wire par_done_reg1180_done;
  wire par_done_reg1181_in;
  wire par_done_reg1181_write_en;
  wire par_done_reg1181_clk;
  wire par_done_reg1181_out;
  wire par_done_reg1181_done;
  wire par_done_reg1182_in;
  wire par_done_reg1182_write_en;
  wire par_done_reg1182_clk;
  wire par_done_reg1182_out;
  wire par_done_reg1182_done;
  wire par_done_reg1183_in;
  wire par_done_reg1183_write_en;
  wire par_done_reg1183_clk;
  wire par_done_reg1183_out;
  wire par_done_reg1183_done;
  wire par_done_reg1184_in;
  wire par_done_reg1184_write_en;
  wire par_done_reg1184_clk;
  wire par_done_reg1184_out;
  wire par_done_reg1184_done;
  wire par_done_reg1185_in;
  wire par_done_reg1185_write_en;
  wire par_done_reg1185_clk;
  wire par_done_reg1185_out;
  wire par_done_reg1185_done;
  wire par_done_reg1186_in;
  wire par_done_reg1186_write_en;
  wire par_done_reg1186_clk;
  wire par_done_reg1186_out;
  wire par_done_reg1186_done;
  wire par_done_reg1187_in;
  wire par_done_reg1187_write_en;
  wire par_done_reg1187_clk;
  wire par_done_reg1187_out;
  wire par_done_reg1187_done;
  wire par_done_reg1188_in;
  wire par_done_reg1188_write_en;
  wire par_done_reg1188_clk;
  wire par_done_reg1188_out;
  wire par_done_reg1188_done;
  wire par_done_reg1189_in;
  wire par_done_reg1189_write_en;
  wire par_done_reg1189_clk;
  wire par_done_reg1189_out;
  wire par_done_reg1189_done;
  wire par_done_reg1190_in;
  wire par_done_reg1190_write_en;
  wire par_done_reg1190_clk;
  wire par_done_reg1190_out;
  wire par_done_reg1190_done;
  wire par_done_reg1191_in;
  wire par_done_reg1191_write_en;
  wire par_done_reg1191_clk;
  wire par_done_reg1191_out;
  wire par_done_reg1191_done;
  wire par_reset28_in;
  wire par_reset28_write_en;
  wire par_reset28_clk;
  wire par_reset28_out;
  wire par_reset28_done;
  wire par_done_reg1192_in;
  wire par_done_reg1192_write_en;
  wire par_done_reg1192_clk;
  wire par_done_reg1192_out;
  wire par_done_reg1192_done;
  wire par_done_reg1193_in;
  wire par_done_reg1193_write_en;
  wire par_done_reg1193_clk;
  wire par_done_reg1193_out;
  wire par_done_reg1193_done;
  wire par_done_reg1194_in;
  wire par_done_reg1194_write_en;
  wire par_done_reg1194_clk;
  wire par_done_reg1194_out;
  wire par_done_reg1194_done;
  wire par_done_reg1195_in;
  wire par_done_reg1195_write_en;
  wire par_done_reg1195_clk;
  wire par_done_reg1195_out;
  wire par_done_reg1195_done;
  wire par_done_reg1196_in;
  wire par_done_reg1196_write_en;
  wire par_done_reg1196_clk;
  wire par_done_reg1196_out;
  wire par_done_reg1196_done;
  wire par_done_reg1197_in;
  wire par_done_reg1197_write_en;
  wire par_done_reg1197_clk;
  wire par_done_reg1197_out;
  wire par_done_reg1197_done;
  wire par_done_reg1198_in;
  wire par_done_reg1198_write_en;
  wire par_done_reg1198_clk;
  wire par_done_reg1198_out;
  wire par_done_reg1198_done;
  wire par_done_reg1199_in;
  wire par_done_reg1199_write_en;
  wire par_done_reg1199_clk;
  wire par_done_reg1199_out;
  wire par_done_reg1199_done;
  wire par_done_reg1200_in;
  wire par_done_reg1200_write_en;
  wire par_done_reg1200_clk;
  wire par_done_reg1200_out;
  wire par_done_reg1200_done;
  wire par_done_reg1201_in;
  wire par_done_reg1201_write_en;
  wire par_done_reg1201_clk;
  wire par_done_reg1201_out;
  wire par_done_reg1201_done;
  wire par_done_reg1202_in;
  wire par_done_reg1202_write_en;
  wire par_done_reg1202_clk;
  wire par_done_reg1202_out;
  wire par_done_reg1202_done;
  wire par_done_reg1203_in;
  wire par_done_reg1203_write_en;
  wire par_done_reg1203_clk;
  wire par_done_reg1203_out;
  wire par_done_reg1203_done;
  wire par_done_reg1204_in;
  wire par_done_reg1204_write_en;
  wire par_done_reg1204_clk;
  wire par_done_reg1204_out;
  wire par_done_reg1204_done;
  wire par_done_reg1205_in;
  wire par_done_reg1205_write_en;
  wire par_done_reg1205_clk;
  wire par_done_reg1205_out;
  wire par_done_reg1205_done;
  wire par_done_reg1206_in;
  wire par_done_reg1206_write_en;
  wire par_done_reg1206_clk;
  wire par_done_reg1206_out;
  wire par_done_reg1206_done;
  wire par_done_reg1207_in;
  wire par_done_reg1207_write_en;
  wire par_done_reg1207_clk;
  wire par_done_reg1207_out;
  wire par_done_reg1207_done;
  wire par_done_reg1208_in;
  wire par_done_reg1208_write_en;
  wire par_done_reg1208_clk;
  wire par_done_reg1208_out;
  wire par_done_reg1208_done;
  wire par_done_reg1209_in;
  wire par_done_reg1209_write_en;
  wire par_done_reg1209_clk;
  wire par_done_reg1209_out;
  wire par_done_reg1209_done;
  wire par_done_reg1210_in;
  wire par_done_reg1210_write_en;
  wire par_done_reg1210_clk;
  wire par_done_reg1210_out;
  wire par_done_reg1210_done;
  wire par_done_reg1211_in;
  wire par_done_reg1211_write_en;
  wire par_done_reg1211_clk;
  wire par_done_reg1211_out;
  wire par_done_reg1211_done;
  wire par_done_reg1212_in;
  wire par_done_reg1212_write_en;
  wire par_done_reg1212_clk;
  wire par_done_reg1212_out;
  wire par_done_reg1212_done;
  wire par_done_reg1213_in;
  wire par_done_reg1213_write_en;
  wire par_done_reg1213_clk;
  wire par_done_reg1213_out;
  wire par_done_reg1213_done;
  wire par_done_reg1214_in;
  wire par_done_reg1214_write_en;
  wire par_done_reg1214_clk;
  wire par_done_reg1214_out;
  wire par_done_reg1214_done;
  wire par_done_reg1215_in;
  wire par_done_reg1215_write_en;
  wire par_done_reg1215_clk;
  wire par_done_reg1215_out;
  wire par_done_reg1215_done;
  wire par_done_reg1216_in;
  wire par_done_reg1216_write_en;
  wire par_done_reg1216_clk;
  wire par_done_reg1216_out;
  wire par_done_reg1216_done;
  wire par_done_reg1217_in;
  wire par_done_reg1217_write_en;
  wire par_done_reg1217_clk;
  wire par_done_reg1217_out;
  wire par_done_reg1217_done;
  wire par_done_reg1218_in;
  wire par_done_reg1218_write_en;
  wire par_done_reg1218_clk;
  wire par_done_reg1218_out;
  wire par_done_reg1218_done;
  wire par_done_reg1219_in;
  wire par_done_reg1219_write_en;
  wire par_done_reg1219_clk;
  wire par_done_reg1219_out;
  wire par_done_reg1219_done;
  wire par_done_reg1220_in;
  wire par_done_reg1220_write_en;
  wire par_done_reg1220_clk;
  wire par_done_reg1220_out;
  wire par_done_reg1220_done;
  wire par_done_reg1221_in;
  wire par_done_reg1221_write_en;
  wire par_done_reg1221_clk;
  wire par_done_reg1221_out;
  wire par_done_reg1221_done;
  wire par_done_reg1222_in;
  wire par_done_reg1222_write_en;
  wire par_done_reg1222_clk;
  wire par_done_reg1222_out;
  wire par_done_reg1222_done;
  wire par_done_reg1223_in;
  wire par_done_reg1223_write_en;
  wire par_done_reg1223_clk;
  wire par_done_reg1223_out;
  wire par_done_reg1223_done;
  wire par_done_reg1224_in;
  wire par_done_reg1224_write_en;
  wire par_done_reg1224_clk;
  wire par_done_reg1224_out;
  wire par_done_reg1224_done;
  wire par_done_reg1225_in;
  wire par_done_reg1225_write_en;
  wire par_done_reg1225_clk;
  wire par_done_reg1225_out;
  wire par_done_reg1225_done;
  wire par_done_reg1226_in;
  wire par_done_reg1226_write_en;
  wire par_done_reg1226_clk;
  wire par_done_reg1226_out;
  wire par_done_reg1226_done;
  wire par_done_reg1227_in;
  wire par_done_reg1227_write_en;
  wire par_done_reg1227_clk;
  wire par_done_reg1227_out;
  wire par_done_reg1227_done;
  wire par_done_reg1228_in;
  wire par_done_reg1228_write_en;
  wire par_done_reg1228_clk;
  wire par_done_reg1228_out;
  wire par_done_reg1228_done;
  wire par_done_reg1229_in;
  wire par_done_reg1229_write_en;
  wire par_done_reg1229_clk;
  wire par_done_reg1229_out;
  wire par_done_reg1229_done;
  wire par_done_reg1230_in;
  wire par_done_reg1230_write_en;
  wire par_done_reg1230_clk;
  wire par_done_reg1230_out;
  wire par_done_reg1230_done;
  wire par_done_reg1231_in;
  wire par_done_reg1231_write_en;
  wire par_done_reg1231_clk;
  wire par_done_reg1231_out;
  wire par_done_reg1231_done;
  wire par_done_reg1232_in;
  wire par_done_reg1232_write_en;
  wire par_done_reg1232_clk;
  wire par_done_reg1232_out;
  wire par_done_reg1232_done;
  wire par_done_reg1233_in;
  wire par_done_reg1233_write_en;
  wire par_done_reg1233_clk;
  wire par_done_reg1233_out;
  wire par_done_reg1233_done;
  wire par_done_reg1234_in;
  wire par_done_reg1234_write_en;
  wire par_done_reg1234_clk;
  wire par_done_reg1234_out;
  wire par_done_reg1234_done;
  wire par_done_reg1235_in;
  wire par_done_reg1235_write_en;
  wire par_done_reg1235_clk;
  wire par_done_reg1235_out;
  wire par_done_reg1235_done;
  wire par_done_reg1236_in;
  wire par_done_reg1236_write_en;
  wire par_done_reg1236_clk;
  wire par_done_reg1236_out;
  wire par_done_reg1236_done;
  wire par_done_reg1237_in;
  wire par_done_reg1237_write_en;
  wire par_done_reg1237_clk;
  wire par_done_reg1237_out;
  wire par_done_reg1237_done;
  wire par_done_reg1238_in;
  wire par_done_reg1238_write_en;
  wire par_done_reg1238_clk;
  wire par_done_reg1238_out;
  wire par_done_reg1238_done;
  wire par_done_reg1239_in;
  wire par_done_reg1239_write_en;
  wire par_done_reg1239_clk;
  wire par_done_reg1239_out;
  wire par_done_reg1239_done;
  wire par_done_reg1240_in;
  wire par_done_reg1240_write_en;
  wire par_done_reg1240_clk;
  wire par_done_reg1240_out;
  wire par_done_reg1240_done;
  wire par_done_reg1241_in;
  wire par_done_reg1241_write_en;
  wire par_done_reg1241_clk;
  wire par_done_reg1241_out;
  wire par_done_reg1241_done;
  wire par_done_reg1242_in;
  wire par_done_reg1242_write_en;
  wire par_done_reg1242_clk;
  wire par_done_reg1242_out;
  wire par_done_reg1242_done;
  wire par_done_reg1243_in;
  wire par_done_reg1243_write_en;
  wire par_done_reg1243_clk;
  wire par_done_reg1243_out;
  wire par_done_reg1243_done;
  wire par_done_reg1244_in;
  wire par_done_reg1244_write_en;
  wire par_done_reg1244_clk;
  wire par_done_reg1244_out;
  wire par_done_reg1244_done;
  wire par_done_reg1245_in;
  wire par_done_reg1245_write_en;
  wire par_done_reg1245_clk;
  wire par_done_reg1245_out;
  wire par_done_reg1245_done;
  wire par_done_reg1246_in;
  wire par_done_reg1246_write_en;
  wire par_done_reg1246_clk;
  wire par_done_reg1246_out;
  wire par_done_reg1246_done;
  wire par_done_reg1247_in;
  wire par_done_reg1247_write_en;
  wire par_done_reg1247_clk;
  wire par_done_reg1247_out;
  wire par_done_reg1247_done;
  wire par_done_reg1248_in;
  wire par_done_reg1248_write_en;
  wire par_done_reg1248_clk;
  wire par_done_reg1248_out;
  wire par_done_reg1248_done;
  wire par_done_reg1249_in;
  wire par_done_reg1249_write_en;
  wire par_done_reg1249_clk;
  wire par_done_reg1249_out;
  wire par_done_reg1249_done;
  wire par_done_reg1250_in;
  wire par_done_reg1250_write_en;
  wire par_done_reg1250_clk;
  wire par_done_reg1250_out;
  wire par_done_reg1250_done;
  wire par_done_reg1251_in;
  wire par_done_reg1251_write_en;
  wire par_done_reg1251_clk;
  wire par_done_reg1251_out;
  wire par_done_reg1251_done;
  wire par_done_reg1252_in;
  wire par_done_reg1252_write_en;
  wire par_done_reg1252_clk;
  wire par_done_reg1252_out;
  wire par_done_reg1252_done;
  wire par_done_reg1253_in;
  wire par_done_reg1253_write_en;
  wire par_done_reg1253_clk;
  wire par_done_reg1253_out;
  wire par_done_reg1253_done;
  wire par_done_reg1254_in;
  wire par_done_reg1254_write_en;
  wire par_done_reg1254_clk;
  wire par_done_reg1254_out;
  wire par_done_reg1254_done;
  wire par_done_reg1255_in;
  wire par_done_reg1255_write_en;
  wire par_done_reg1255_clk;
  wire par_done_reg1255_out;
  wire par_done_reg1255_done;
  wire par_done_reg1256_in;
  wire par_done_reg1256_write_en;
  wire par_done_reg1256_clk;
  wire par_done_reg1256_out;
  wire par_done_reg1256_done;
  wire par_done_reg1257_in;
  wire par_done_reg1257_write_en;
  wire par_done_reg1257_clk;
  wire par_done_reg1257_out;
  wire par_done_reg1257_done;
  wire par_done_reg1258_in;
  wire par_done_reg1258_write_en;
  wire par_done_reg1258_clk;
  wire par_done_reg1258_out;
  wire par_done_reg1258_done;
  wire par_done_reg1259_in;
  wire par_done_reg1259_write_en;
  wire par_done_reg1259_clk;
  wire par_done_reg1259_out;
  wire par_done_reg1259_done;
  wire par_done_reg1260_in;
  wire par_done_reg1260_write_en;
  wire par_done_reg1260_clk;
  wire par_done_reg1260_out;
  wire par_done_reg1260_done;
  wire par_done_reg1261_in;
  wire par_done_reg1261_write_en;
  wire par_done_reg1261_clk;
  wire par_done_reg1261_out;
  wire par_done_reg1261_done;
  wire par_done_reg1262_in;
  wire par_done_reg1262_write_en;
  wire par_done_reg1262_clk;
  wire par_done_reg1262_out;
  wire par_done_reg1262_done;
  wire par_done_reg1263_in;
  wire par_done_reg1263_write_en;
  wire par_done_reg1263_clk;
  wire par_done_reg1263_out;
  wire par_done_reg1263_done;
  wire par_done_reg1264_in;
  wire par_done_reg1264_write_en;
  wire par_done_reg1264_clk;
  wire par_done_reg1264_out;
  wire par_done_reg1264_done;
  wire par_done_reg1265_in;
  wire par_done_reg1265_write_en;
  wire par_done_reg1265_clk;
  wire par_done_reg1265_out;
  wire par_done_reg1265_done;
  wire par_done_reg1266_in;
  wire par_done_reg1266_write_en;
  wire par_done_reg1266_clk;
  wire par_done_reg1266_out;
  wire par_done_reg1266_done;
  wire par_done_reg1267_in;
  wire par_done_reg1267_write_en;
  wire par_done_reg1267_clk;
  wire par_done_reg1267_out;
  wire par_done_reg1267_done;
  wire par_done_reg1268_in;
  wire par_done_reg1268_write_en;
  wire par_done_reg1268_clk;
  wire par_done_reg1268_out;
  wire par_done_reg1268_done;
  wire par_done_reg1269_in;
  wire par_done_reg1269_write_en;
  wire par_done_reg1269_clk;
  wire par_done_reg1269_out;
  wire par_done_reg1269_done;
  wire par_done_reg1270_in;
  wire par_done_reg1270_write_en;
  wire par_done_reg1270_clk;
  wire par_done_reg1270_out;
  wire par_done_reg1270_done;
  wire par_done_reg1271_in;
  wire par_done_reg1271_write_en;
  wire par_done_reg1271_clk;
  wire par_done_reg1271_out;
  wire par_done_reg1271_done;
  wire par_done_reg1272_in;
  wire par_done_reg1272_write_en;
  wire par_done_reg1272_clk;
  wire par_done_reg1272_out;
  wire par_done_reg1272_done;
  wire par_done_reg1273_in;
  wire par_done_reg1273_write_en;
  wire par_done_reg1273_clk;
  wire par_done_reg1273_out;
  wire par_done_reg1273_done;
  wire par_done_reg1274_in;
  wire par_done_reg1274_write_en;
  wire par_done_reg1274_clk;
  wire par_done_reg1274_out;
  wire par_done_reg1274_done;
  wire par_done_reg1275_in;
  wire par_done_reg1275_write_en;
  wire par_done_reg1275_clk;
  wire par_done_reg1275_out;
  wire par_done_reg1275_done;
  wire par_reset29_in;
  wire par_reset29_write_en;
  wire par_reset29_clk;
  wire par_reset29_out;
  wire par_reset29_done;
  wire par_done_reg1276_in;
  wire par_done_reg1276_write_en;
  wire par_done_reg1276_clk;
  wire par_done_reg1276_out;
  wire par_done_reg1276_done;
  wire par_done_reg1277_in;
  wire par_done_reg1277_write_en;
  wire par_done_reg1277_clk;
  wire par_done_reg1277_out;
  wire par_done_reg1277_done;
  wire par_done_reg1278_in;
  wire par_done_reg1278_write_en;
  wire par_done_reg1278_clk;
  wire par_done_reg1278_out;
  wire par_done_reg1278_done;
  wire par_done_reg1279_in;
  wire par_done_reg1279_write_en;
  wire par_done_reg1279_clk;
  wire par_done_reg1279_out;
  wire par_done_reg1279_done;
  wire par_done_reg1280_in;
  wire par_done_reg1280_write_en;
  wire par_done_reg1280_clk;
  wire par_done_reg1280_out;
  wire par_done_reg1280_done;
  wire par_done_reg1281_in;
  wire par_done_reg1281_write_en;
  wire par_done_reg1281_clk;
  wire par_done_reg1281_out;
  wire par_done_reg1281_done;
  wire par_done_reg1282_in;
  wire par_done_reg1282_write_en;
  wire par_done_reg1282_clk;
  wire par_done_reg1282_out;
  wire par_done_reg1282_done;
  wire par_done_reg1283_in;
  wire par_done_reg1283_write_en;
  wire par_done_reg1283_clk;
  wire par_done_reg1283_out;
  wire par_done_reg1283_done;
  wire par_done_reg1284_in;
  wire par_done_reg1284_write_en;
  wire par_done_reg1284_clk;
  wire par_done_reg1284_out;
  wire par_done_reg1284_done;
  wire par_done_reg1285_in;
  wire par_done_reg1285_write_en;
  wire par_done_reg1285_clk;
  wire par_done_reg1285_out;
  wire par_done_reg1285_done;
  wire par_done_reg1286_in;
  wire par_done_reg1286_write_en;
  wire par_done_reg1286_clk;
  wire par_done_reg1286_out;
  wire par_done_reg1286_done;
  wire par_done_reg1287_in;
  wire par_done_reg1287_write_en;
  wire par_done_reg1287_clk;
  wire par_done_reg1287_out;
  wire par_done_reg1287_done;
  wire par_done_reg1288_in;
  wire par_done_reg1288_write_en;
  wire par_done_reg1288_clk;
  wire par_done_reg1288_out;
  wire par_done_reg1288_done;
  wire par_done_reg1289_in;
  wire par_done_reg1289_write_en;
  wire par_done_reg1289_clk;
  wire par_done_reg1289_out;
  wire par_done_reg1289_done;
  wire par_done_reg1290_in;
  wire par_done_reg1290_write_en;
  wire par_done_reg1290_clk;
  wire par_done_reg1290_out;
  wire par_done_reg1290_done;
  wire par_done_reg1291_in;
  wire par_done_reg1291_write_en;
  wire par_done_reg1291_clk;
  wire par_done_reg1291_out;
  wire par_done_reg1291_done;
  wire par_done_reg1292_in;
  wire par_done_reg1292_write_en;
  wire par_done_reg1292_clk;
  wire par_done_reg1292_out;
  wire par_done_reg1292_done;
  wire par_done_reg1293_in;
  wire par_done_reg1293_write_en;
  wire par_done_reg1293_clk;
  wire par_done_reg1293_out;
  wire par_done_reg1293_done;
  wire par_done_reg1294_in;
  wire par_done_reg1294_write_en;
  wire par_done_reg1294_clk;
  wire par_done_reg1294_out;
  wire par_done_reg1294_done;
  wire par_done_reg1295_in;
  wire par_done_reg1295_write_en;
  wire par_done_reg1295_clk;
  wire par_done_reg1295_out;
  wire par_done_reg1295_done;
  wire par_done_reg1296_in;
  wire par_done_reg1296_write_en;
  wire par_done_reg1296_clk;
  wire par_done_reg1296_out;
  wire par_done_reg1296_done;
  wire par_done_reg1297_in;
  wire par_done_reg1297_write_en;
  wire par_done_reg1297_clk;
  wire par_done_reg1297_out;
  wire par_done_reg1297_done;
  wire par_done_reg1298_in;
  wire par_done_reg1298_write_en;
  wire par_done_reg1298_clk;
  wire par_done_reg1298_out;
  wire par_done_reg1298_done;
  wire par_done_reg1299_in;
  wire par_done_reg1299_write_en;
  wire par_done_reg1299_clk;
  wire par_done_reg1299_out;
  wire par_done_reg1299_done;
  wire par_done_reg1300_in;
  wire par_done_reg1300_write_en;
  wire par_done_reg1300_clk;
  wire par_done_reg1300_out;
  wire par_done_reg1300_done;
  wire par_done_reg1301_in;
  wire par_done_reg1301_write_en;
  wire par_done_reg1301_clk;
  wire par_done_reg1301_out;
  wire par_done_reg1301_done;
  wire par_done_reg1302_in;
  wire par_done_reg1302_write_en;
  wire par_done_reg1302_clk;
  wire par_done_reg1302_out;
  wire par_done_reg1302_done;
  wire par_done_reg1303_in;
  wire par_done_reg1303_write_en;
  wire par_done_reg1303_clk;
  wire par_done_reg1303_out;
  wire par_done_reg1303_done;
  wire par_done_reg1304_in;
  wire par_done_reg1304_write_en;
  wire par_done_reg1304_clk;
  wire par_done_reg1304_out;
  wire par_done_reg1304_done;
  wire par_done_reg1305_in;
  wire par_done_reg1305_write_en;
  wire par_done_reg1305_clk;
  wire par_done_reg1305_out;
  wire par_done_reg1305_done;
  wire par_done_reg1306_in;
  wire par_done_reg1306_write_en;
  wire par_done_reg1306_clk;
  wire par_done_reg1306_out;
  wire par_done_reg1306_done;
  wire par_done_reg1307_in;
  wire par_done_reg1307_write_en;
  wire par_done_reg1307_clk;
  wire par_done_reg1307_out;
  wire par_done_reg1307_done;
  wire par_done_reg1308_in;
  wire par_done_reg1308_write_en;
  wire par_done_reg1308_clk;
  wire par_done_reg1308_out;
  wire par_done_reg1308_done;
  wire par_done_reg1309_in;
  wire par_done_reg1309_write_en;
  wire par_done_reg1309_clk;
  wire par_done_reg1309_out;
  wire par_done_reg1309_done;
  wire par_done_reg1310_in;
  wire par_done_reg1310_write_en;
  wire par_done_reg1310_clk;
  wire par_done_reg1310_out;
  wire par_done_reg1310_done;
  wire par_done_reg1311_in;
  wire par_done_reg1311_write_en;
  wire par_done_reg1311_clk;
  wire par_done_reg1311_out;
  wire par_done_reg1311_done;
  wire par_done_reg1312_in;
  wire par_done_reg1312_write_en;
  wire par_done_reg1312_clk;
  wire par_done_reg1312_out;
  wire par_done_reg1312_done;
  wire par_done_reg1313_in;
  wire par_done_reg1313_write_en;
  wire par_done_reg1313_clk;
  wire par_done_reg1313_out;
  wire par_done_reg1313_done;
  wire par_done_reg1314_in;
  wire par_done_reg1314_write_en;
  wire par_done_reg1314_clk;
  wire par_done_reg1314_out;
  wire par_done_reg1314_done;
  wire par_done_reg1315_in;
  wire par_done_reg1315_write_en;
  wire par_done_reg1315_clk;
  wire par_done_reg1315_out;
  wire par_done_reg1315_done;
  wire par_done_reg1316_in;
  wire par_done_reg1316_write_en;
  wire par_done_reg1316_clk;
  wire par_done_reg1316_out;
  wire par_done_reg1316_done;
  wire par_done_reg1317_in;
  wire par_done_reg1317_write_en;
  wire par_done_reg1317_clk;
  wire par_done_reg1317_out;
  wire par_done_reg1317_done;
  wire par_done_reg1318_in;
  wire par_done_reg1318_write_en;
  wire par_done_reg1318_clk;
  wire par_done_reg1318_out;
  wire par_done_reg1318_done;
  wire par_done_reg1319_in;
  wire par_done_reg1319_write_en;
  wire par_done_reg1319_clk;
  wire par_done_reg1319_out;
  wire par_done_reg1319_done;
  wire par_reset30_in;
  wire par_reset30_write_en;
  wire par_reset30_clk;
  wire par_reset30_out;
  wire par_reset30_done;
  wire par_done_reg1320_in;
  wire par_done_reg1320_write_en;
  wire par_done_reg1320_clk;
  wire par_done_reg1320_out;
  wire par_done_reg1320_done;
  wire par_done_reg1321_in;
  wire par_done_reg1321_write_en;
  wire par_done_reg1321_clk;
  wire par_done_reg1321_out;
  wire par_done_reg1321_done;
  wire par_done_reg1322_in;
  wire par_done_reg1322_write_en;
  wire par_done_reg1322_clk;
  wire par_done_reg1322_out;
  wire par_done_reg1322_done;
  wire par_done_reg1323_in;
  wire par_done_reg1323_write_en;
  wire par_done_reg1323_clk;
  wire par_done_reg1323_out;
  wire par_done_reg1323_done;
  wire par_done_reg1324_in;
  wire par_done_reg1324_write_en;
  wire par_done_reg1324_clk;
  wire par_done_reg1324_out;
  wire par_done_reg1324_done;
  wire par_done_reg1325_in;
  wire par_done_reg1325_write_en;
  wire par_done_reg1325_clk;
  wire par_done_reg1325_out;
  wire par_done_reg1325_done;
  wire par_done_reg1326_in;
  wire par_done_reg1326_write_en;
  wire par_done_reg1326_clk;
  wire par_done_reg1326_out;
  wire par_done_reg1326_done;
  wire par_done_reg1327_in;
  wire par_done_reg1327_write_en;
  wire par_done_reg1327_clk;
  wire par_done_reg1327_out;
  wire par_done_reg1327_done;
  wire par_done_reg1328_in;
  wire par_done_reg1328_write_en;
  wire par_done_reg1328_clk;
  wire par_done_reg1328_out;
  wire par_done_reg1328_done;
  wire par_done_reg1329_in;
  wire par_done_reg1329_write_en;
  wire par_done_reg1329_clk;
  wire par_done_reg1329_out;
  wire par_done_reg1329_done;
  wire par_done_reg1330_in;
  wire par_done_reg1330_write_en;
  wire par_done_reg1330_clk;
  wire par_done_reg1330_out;
  wire par_done_reg1330_done;
  wire par_done_reg1331_in;
  wire par_done_reg1331_write_en;
  wire par_done_reg1331_clk;
  wire par_done_reg1331_out;
  wire par_done_reg1331_done;
  wire par_done_reg1332_in;
  wire par_done_reg1332_write_en;
  wire par_done_reg1332_clk;
  wire par_done_reg1332_out;
  wire par_done_reg1332_done;
  wire par_done_reg1333_in;
  wire par_done_reg1333_write_en;
  wire par_done_reg1333_clk;
  wire par_done_reg1333_out;
  wire par_done_reg1333_done;
  wire par_done_reg1334_in;
  wire par_done_reg1334_write_en;
  wire par_done_reg1334_clk;
  wire par_done_reg1334_out;
  wire par_done_reg1334_done;
  wire par_done_reg1335_in;
  wire par_done_reg1335_write_en;
  wire par_done_reg1335_clk;
  wire par_done_reg1335_out;
  wire par_done_reg1335_done;
  wire par_done_reg1336_in;
  wire par_done_reg1336_write_en;
  wire par_done_reg1336_clk;
  wire par_done_reg1336_out;
  wire par_done_reg1336_done;
  wire par_done_reg1337_in;
  wire par_done_reg1337_write_en;
  wire par_done_reg1337_clk;
  wire par_done_reg1337_out;
  wire par_done_reg1337_done;
  wire par_done_reg1338_in;
  wire par_done_reg1338_write_en;
  wire par_done_reg1338_clk;
  wire par_done_reg1338_out;
  wire par_done_reg1338_done;
  wire par_done_reg1339_in;
  wire par_done_reg1339_write_en;
  wire par_done_reg1339_clk;
  wire par_done_reg1339_out;
  wire par_done_reg1339_done;
  wire par_done_reg1340_in;
  wire par_done_reg1340_write_en;
  wire par_done_reg1340_clk;
  wire par_done_reg1340_out;
  wire par_done_reg1340_done;
  wire par_done_reg1341_in;
  wire par_done_reg1341_write_en;
  wire par_done_reg1341_clk;
  wire par_done_reg1341_out;
  wire par_done_reg1341_done;
  wire par_done_reg1342_in;
  wire par_done_reg1342_write_en;
  wire par_done_reg1342_clk;
  wire par_done_reg1342_out;
  wire par_done_reg1342_done;
  wire par_done_reg1343_in;
  wire par_done_reg1343_write_en;
  wire par_done_reg1343_clk;
  wire par_done_reg1343_out;
  wire par_done_reg1343_done;
  wire par_done_reg1344_in;
  wire par_done_reg1344_write_en;
  wire par_done_reg1344_clk;
  wire par_done_reg1344_out;
  wire par_done_reg1344_done;
  wire par_done_reg1345_in;
  wire par_done_reg1345_write_en;
  wire par_done_reg1345_clk;
  wire par_done_reg1345_out;
  wire par_done_reg1345_done;
  wire par_done_reg1346_in;
  wire par_done_reg1346_write_en;
  wire par_done_reg1346_clk;
  wire par_done_reg1346_out;
  wire par_done_reg1346_done;
  wire par_done_reg1347_in;
  wire par_done_reg1347_write_en;
  wire par_done_reg1347_clk;
  wire par_done_reg1347_out;
  wire par_done_reg1347_done;
  wire par_done_reg1348_in;
  wire par_done_reg1348_write_en;
  wire par_done_reg1348_clk;
  wire par_done_reg1348_out;
  wire par_done_reg1348_done;
  wire par_done_reg1349_in;
  wire par_done_reg1349_write_en;
  wire par_done_reg1349_clk;
  wire par_done_reg1349_out;
  wire par_done_reg1349_done;
  wire par_done_reg1350_in;
  wire par_done_reg1350_write_en;
  wire par_done_reg1350_clk;
  wire par_done_reg1350_out;
  wire par_done_reg1350_done;
  wire par_done_reg1351_in;
  wire par_done_reg1351_write_en;
  wire par_done_reg1351_clk;
  wire par_done_reg1351_out;
  wire par_done_reg1351_done;
  wire par_done_reg1352_in;
  wire par_done_reg1352_write_en;
  wire par_done_reg1352_clk;
  wire par_done_reg1352_out;
  wire par_done_reg1352_done;
  wire par_done_reg1353_in;
  wire par_done_reg1353_write_en;
  wire par_done_reg1353_clk;
  wire par_done_reg1353_out;
  wire par_done_reg1353_done;
  wire par_done_reg1354_in;
  wire par_done_reg1354_write_en;
  wire par_done_reg1354_clk;
  wire par_done_reg1354_out;
  wire par_done_reg1354_done;
  wire par_done_reg1355_in;
  wire par_done_reg1355_write_en;
  wire par_done_reg1355_clk;
  wire par_done_reg1355_out;
  wire par_done_reg1355_done;
  wire par_done_reg1356_in;
  wire par_done_reg1356_write_en;
  wire par_done_reg1356_clk;
  wire par_done_reg1356_out;
  wire par_done_reg1356_done;
  wire par_done_reg1357_in;
  wire par_done_reg1357_write_en;
  wire par_done_reg1357_clk;
  wire par_done_reg1357_out;
  wire par_done_reg1357_done;
  wire par_done_reg1358_in;
  wire par_done_reg1358_write_en;
  wire par_done_reg1358_clk;
  wire par_done_reg1358_out;
  wire par_done_reg1358_done;
  wire par_done_reg1359_in;
  wire par_done_reg1359_write_en;
  wire par_done_reg1359_clk;
  wire par_done_reg1359_out;
  wire par_done_reg1359_done;
  wire par_done_reg1360_in;
  wire par_done_reg1360_write_en;
  wire par_done_reg1360_clk;
  wire par_done_reg1360_out;
  wire par_done_reg1360_done;
  wire par_done_reg1361_in;
  wire par_done_reg1361_write_en;
  wire par_done_reg1361_clk;
  wire par_done_reg1361_out;
  wire par_done_reg1361_done;
  wire par_done_reg1362_in;
  wire par_done_reg1362_write_en;
  wire par_done_reg1362_clk;
  wire par_done_reg1362_out;
  wire par_done_reg1362_done;
  wire par_done_reg1363_in;
  wire par_done_reg1363_write_en;
  wire par_done_reg1363_clk;
  wire par_done_reg1363_out;
  wire par_done_reg1363_done;
  wire par_done_reg1364_in;
  wire par_done_reg1364_write_en;
  wire par_done_reg1364_clk;
  wire par_done_reg1364_out;
  wire par_done_reg1364_done;
  wire par_done_reg1365_in;
  wire par_done_reg1365_write_en;
  wire par_done_reg1365_clk;
  wire par_done_reg1365_out;
  wire par_done_reg1365_done;
  wire par_done_reg1366_in;
  wire par_done_reg1366_write_en;
  wire par_done_reg1366_clk;
  wire par_done_reg1366_out;
  wire par_done_reg1366_done;
  wire par_done_reg1367_in;
  wire par_done_reg1367_write_en;
  wire par_done_reg1367_clk;
  wire par_done_reg1367_out;
  wire par_done_reg1367_done;
  wire par_done_reg1368_in;
  wire par_done_reg1368_write_en;
  wire par_done_reg1368_clk;
  wire par_done_reg1368_out;
  wire par_done_reg1368_done;
  wire par_done_reg1369_in;
  wire par_done_reg1369_write_en;
  wire par_done_reg1369_clk;
  wire par_done_reg1369_out;
  wire par_done_reg1369_done;
  wire par_done_reg1370_in;
  wire par_done_reg1370_write_en;
  wire par_done_reg1370_clk;
  wire par_done_reg1370_out;
  wire par_done_reg1370_done;
  wire par_done_reg1371_in;
  wire par_done_reg1371_write_en;
  wire par_done_reg1371_clk;
  wire par_done_reg1371_out;
  wire par_done_reg1371_done;
  wire par_done_reg1372_in;
  wire par_done_reg1372_write_en;
  wire par_done_reg1372_clk;
  wire par_done_reg1372_out;
  wire par_done_reg1372_done;
  wire par_done_reg1373_in;
  wire par_done_reg1373_write_en;
  wire par_done_reg1373_clk;
  wire par_done_reg1373_out;
  wire par_done_reg1373_done;
  wire par_done_reg1374_in;
  wire par_done_reg1374_write_en;
  wire par_done_reg1374_clk;
  wire par_done_reg1374_out;
  wire par_done_reg1374_done;
  wire par_done_reg1375_in;
  wire par_done_reg1375_write_en;
  wire par_done_reg1375_clk;
  wire par_done_reg1375_out;
  wire par_done_reg1375_done;
  wire par_done_reg1376_in;
  wire par_done_reg1376_write_en;
  wire par_done_reg1376_clk;
  wire par_done_reg1376_out;
  wire par_done_reg1376_done;
  wire par_done_reg1377_in;
  wire par_done_reg1377_write_en;
  wire par_done_reg1377_clk;
  wire par_done_reg1377_out;
  wire par_done_reg1377_done;
  wire par_done_reg1378_in;
  wire par_done_reg1378_write_en;
  wire par_done_reg1378_clk;
  wire par_done_reg1378_out;
  wire par_done_reg1378_done;
  wire par_done_reg1379_in;
  wire par_done_reg1379_write_en;
  wire par_done_reg1379_clk;
  wire par_done_reg1379_out;
  wire par_done_reg1379_done;
  wire par_done_reg1380_in;
  wire par_done_reg1380_write_en;
  wire par_done_reg1380_clk;
  wire par_done_reg1380_out;
  wire par_done_reg1380_done;
  wire par_done_reg1381_in;
  wire par_done_reg1381_write_en;
  wire par_done_reg1381_clk;
  wire par_done_reg1381_out;
  wire par_done_reg1381_done;
  wire par_done_reg1382_in;
  wire par_done_reg1382_write_en;
  wire par_done_reg1382_clk;
  wire par_done_reg1382_out;
  wire par_done_reg1382_done;
  wire par_done_reg1383_in;
  wire par_done_reg1383_write_en;
  wire par_done_reg1383_clk;
  wire par_done_reg1383_out;
  wire par_done_reg1383_done;
  wire par_done_reg1384_in;
  wire par_done_reg1384_write_en;
  wire par_done_reg1384_clk;
  wire par_done_reg1384_out;
  wire par_done_reg1384_done;
  wire par_done_reg1385_in;
  wire par_done_reg1385_write_en;
  wire par_done_reg1385_clk;
  wire par_done_reg1385_out;
  wire par_done_reg1385_done;
  wire par_done_reg1386_in;
  wire par_done_reg1386_write_en;
  wire par_done_reg1386_clk;
  wire par_done_reg1386_out;
  wire par_done_reg1386_done;
  wire par_done_reg1387_in;
  wire par_done_reg1387_write_en;
  wire par_done_reg1387_clk;
  wire par_done_reg1387_out;
  wire par_done_reg1387_done;
  wire par_done_reg1388_in;
  wire par_done_reg1388_write_en;
  wire par_done_reg1388_clk;
  wire par_done_reg1388_out;
  wire par_done_reg1388_done;
  wire par_done_reg1389_in;
  wire par_done_reg1389_write_en;
  wire par_done_reg1389_clk;
  wire par_done_reg1389_out;
  wire par_done_reg1389_done;
  wire par_done_reg1390_in;
  wire par_done_reg1390_write_en;
  wire par_done_reg1390_clk;
  wire par_done_reg1390_out;
  wire par_done_reg1390_done;
  wire par_done_reg1391_in;
  wire par_done_reg1391_write_en;
  wire par_done_reg1391_clk;
  wire par_done_reg1391_out;
  wire par_done_reg1391_done;
  wire par_reset31_in;
  wire par_reset31_write_en;
  wire par_reset31_clk;
  wire par_reset31_out;
  wire par_reset31_done;
  wire par_done_reg1392_in;
  wire par_done_reg1392_write_en;
  wire par_done_reg1392_clk;
  wire par_done_reg1392_out;
  wire par_done_reg1392_done;
  wire par_done_reg1393_in;
  wire par_done_reg1393_write_en;
  wire par_done_reg1393_clk;
  wire par_done_reg1393_out;
  wire par_done_reg1393_done;
  wire par_done_reg1394_in;
  wire par_done_reg1394_write_en;
  wire par_done_reg1394_clk;
  wire par_done_reg1394_out;
  wire par_done_reg1394_done;
  wire par_done_reg1395_in;
  wire par_done_reg1395_write_en;
  wire par_done_reg1395_clk;
  wire par_done_reg1395_out;
  wire par_done_reg1395_done;
  wire par_done_reg1396_in;
  wire par_done_reg1396_write_en;
  wire par_done_reg1396_clk;
  wire par_done_reg1396_out;
  wire par_done_reg1396_done;
  wire par_done_reg1397_in;
  wire par_done_reg1397_write_en;
  wire par_done_reg1397_clk;
  wire par_done_reg1397_out;
  wire par_done_reg1397_done;
  wire par_done_reg1398_in;
  wire par_done_reg1398_write_en;
  wire par_done_reg1398_clk;
  wire par_done_reg1398_out;
  wire par_done_reg1398_done;
  wire par_done_reg1399_in;
  wire par_done_reg1399_write_en;
  wire par_done_reg1399_clk;
  wire par_done_reg1399_out;
  wire par_done_reg1399_done;
  wire par_done_reg1400_in;
  wire par_done_reg1400_write_en;
  wire par_done_reg1400_clk;
  wire par_done_reg1400_out;
  wire par_done_reg1400_done;
  wire par_done_reg1401_in;
  wire par_done_reg1401_write_en;
  wire par_done_reg1401_clk;
  wire par_done_reg1401_out;
  wire par_done_reg1401_done;
  wire par_done_reg1402_in;
  wire par_done_reg1402_write_en;
  wire par_done_reg1402_clk;
  wire par_done_reg1402_out;
  wire par_done_reg1402_done;
  wire par_done_reg1403_in;
  wire par_done_reg1403_write_en;
  wire par_done_reg1403_clk;
  wire par_done_reg1403_out;
  wire par_done_reg1403_done;
  wire par_done_reg1404_in;
  wire par_done_reg1404_write_en;
  wire par_done_reg1404_clk;
  wire par_done_reg1404_out;
  wire par_done_reg1404_done;
  wire par_done_reg1405_in;
  wire par_done_reg1405_write_en;
  wire par_done_reg1405_clk;
  wire par_done_reg1405_out;
  wire par_done_reg1405_done;
  wire par_done_reg1406_in;
  wire par_done_reg1406_write_en;
  wire par_done_reg1406_clk;
  wire par_done_reg1406_out;
  wire par_done_reg1406_done;
  wire par_done_reg1407_in;
  wire par_done_reg1407_write_en;
  wire par_done_reg1407_clk;
  wire par_done_reg1407_out;
  wire par_done_reg1407_done;
  wire par_done_reg1408_in;
  wire par_done_reg1408_write_en;
  wire par_done_reg1408_clk;
  wire par_done_reg1408_out;
  wire par_done_reg1408_done;
  wire par_done_reg1409_in;
  wire par_done_reg1409_write_en;
  wire par_done_reg1409_clk;
  wire par_done_reg1409_out;
  wire par_done_reg1409_done;
  wire par_done_reg1410_in;
  wire par_done_reg1410_write_en;
  wire par_done_reg1410_clk;
  wire par_done_reg1410_out;
  wire par_done_reg1410_done;
  wire par_done_reg1411_in;
  wire par_done_reg1411_write_en;
  wire par_done_reg1411_clk;
  wire par_done_reg1411_out;
  wire par_done_reg1411_done;
  wire par_done_reg1412_in;
  wire par_done_reg1412_write_en;
  wire par_done_reg1412_clk;
  wire par_done_reg1412_out;
  wire par_done_reg1412_done;
  wire par_done_reg1413_in;
  wire par_done_reg1413_write_en;
  wire par_done_reg1413_clk;
  wire par_done_reg1413_out;
  wire par_done_reg1413_done;
  wire par_done_reg1414_in;
  wire par_done_reg1414_write_en;
  wire par_done_reg1414_clk;
  wire par_done_reg1414_out;
  wire par_done_reg1414_done;
  wire par_done_reg1415_in;
  wire par_done_reg1415_write_en;
  wire par_done_reg1415_clk;
  wire par_done_reg1415_out;
  wire par_done_reg1415_done;
  wire par_done_reg1416_in;
  wire par_done_reg1416_write_en;
  wire par_done_reg1416_clk;
  wire par_done_reg1416_out;
  wire par_done_reg1416_done;
  wire par_done_reg1417_in;
  wire par_done_reg1417_write_en;
  wire par_done_reg1417_clk;
  wire par_done_reg1417_out;
  wire par_done_reg1417_done;
  wire par_done_reg1418_in;
  wire par_done_reg1418_write_en;
  wire par_done_reg1418_clk;
  wire par_done_reg1418_out;
  wire par_done_reg1418_done;
  wire par_done_reg1419_in;
  wire par_done_reg1419_write_en;
  wire par_done_reg1419_clk;
  wire par_done_reg1419_out;
  wire par_done_reg1419_done;
  wire par_done_reg1420_in;
  wire par_done_reg1420_write_en;
  wire par_done_reg1420_clk;
  wire par_done_reg1420_out;
  wire par_done_reg1420_done;
  wire par_done_reg1421_in;
  wire par_done_reg1421_write_en;
  wire par_done_reg1421_clk;
  wire par_done_reg1421_out;
  wire par_done_reg1421_done;
  wire par_done_reg1422_in;
  wire par_done_reg1422_write_en;
  wire par_done_reg1422_clk;
  wire par_done_reg1422_out;
  wire par_done_reg1422_done;
  wire par_done_reg1423_in;
  wire par_done_reg1423_write_en;
  wire par_done_reg1423_clk;
  wire par_done_reg1423_out;
  wire par_done_reg1423_done;
  wire par_done_reg1424_in;
  wire par_done_reg1424_write_en;
  wire par_done_reg1424_clk;
  wire par_done_reg1424_out;
  wire par_done_reg1424_done;
  wire par_done_reg1425_in;
  wire par_done_reg1425_write_en;
  wire par_done_reg1425_clk;
  wire par_done_reg1425_out;
  wire par_done_reg1425_done;
  wire par_done_reg1426_in;
  wire par_done_reg1426_write_en;
  wire par_done_reg1426_clk;
  wire par_done_reg1426_out;
  wire par_done_reg1426_done;
  wire par_done_reg1427_in;
  wire par_done_reg1427_write_en;
  wire par_done_reg1427_clk;
  wire par_done_reg1427_out;
  wire par_done_reg1427_done;
  wire par_reset32_in;
  wire par_reset32_write_en;
  wire par_reset32_clk;
  wire par_reset32_out;
  wire par_reset32_done;
  wire par_done_reg1428_in;
  wire par_done_reg1428_write_en;
  wire par_done_reg1428_clk;
  wire par_done_reg1428_out;
  wire par_done_reg1428_done;
  wire par_done_reg1429_in;
  wire par_done_reg1429_write_en;
  wire par_done_reg1429_clk;
  wire par_done_reg1429_out;
  wire par_done_reg1429_done;
  wire par_done_reg1430_in;
  wire par_done_reg1430_write_en;
  wire par_done_reg1430_clk;
  wire par_done_reg1430_out;
  wire par_done_reg1430_done;
  wire par_done_reg1431_in;
  wire par_done_reg1431_write_en;
  wire par_done_reg1431_clk;
  wire par_done_reg1431_out;
  wire par_done_reg1431_done;
  wire par_done_reg1432_in;
  wire par_done_reg1432_write_en;
  wire par_done_reg1432_clk;
  wire par_done_reg1432_out;
  wire par_done_reg1432_done;
  wire par_done_reg1433_in;
  wire par_done_reg1433_write_en;
  wire par_done_reg1433_clk;
  wire par_done_reg1433_out;
  wire par_done_reg1433_done;
  wire par_done_reg1434_in;
  wire par_done_reg1434_write_en;
  wire par_done_reg1434_clk;
  wire par_done_reg1434_out;
  wire par_done_reg1434_done;
  wire par_done_reg1435_in;
  wire par_done_reg1435_write_en;
  wire par_done_reg1435_clk;
  wire par_done_reg1435_out;
  wire par_done_reg1435_done;
  wire par_done_reg1436_in;
  wire par_done_reg1436_write_en;
  wire par_done_reg1436_clk;
  wire par_done_reg1436_out;
  wire par_done_reg1436_done;
  wire par_done_reg1437_in;
  wire par_done_reg1437_write_en;
  wire par_done_reg1437_clk;
  wire par_done_reg1437_out;
  wire par_done_reg1437_done;
  wire par_done_reg1438_in;
  wire par_done_reg1438_write_en;
  wire par_done_reg1438_clk;
  wire par_done_reg1438_out;
  wire par_done_reg1438_done;
  wire par_done_reg1439_in;
  wire par_done_reg1439_write_en;
  wire par_done_reg1439_clk;
  wire par_done_reg1439_out;
  wire par_done_reg1439_done;
  wire par_done_reg1440_in;
  wire par_done_reg1440_write_en;
  wire par_done_reg1440_clk;
  wire par_done_reg1440_out;
  wire par_done_reg1440_done;
  wire par_done_reg1441_in;
  wire par_done_reg1441_write_en;
  wire par_done_reg1441_clk;
  wire par_done_reg1441_out;
  wire par_done_reg1441_done;
  wire par_done_reg1442_in;
  wire par_done_reg1442_write_en;
  wire par_done_reg1442_clk;
  wire par_done_reg1442_out;
  wire par_done_reg1442_done;
  wire par_done_reg1443_in;
  wire par_done_reg1443_write_en;
  wire par_done_reg1443_clk;
  wire par_done_reg1443_out;
  wire par_done_reg1443_done;
  wire par_done_reg1444_in;
  wire par_done_reg1444_write_en;
  wire par_done_reg1444_clk;
  wire par_done_reg1444_out;
  wire par_done_reg1444_done;
  wire par_done_reg1445_in;
  wire par_done_reg1445_write_en;
  wire par_done_reg1445_clk;
  wire par_done_reg1445_out;
  wire par_done_reg1445_done;
  wire par_done_reg1446_in;
  wire par_done_reg1446_write_en;
  wire par_done_reg1446_clk;
  wire par_done_reg1446_out;
  wire par_done_reg1446_done;
  wire par_done_reg1447_in;
  wire par_done_reg1447_write_en;
  wire par_done_reg1447_clk;
  wire par_done_reg1447_out;
  wire par_done_reg1447_done;
  wire par_done_reg1448_in;
  wire par_done_reg1448_write_en;
  wire par_done_reg1448_clk;
  wire par_done_reg1448_out;
  wire par_done_reg1448_done;
  wire par_done_reg1449_in;
  wire par_done_reg1449_write_en;
  wire par_done_reg1449_clk;
  wire par_done_reg1449_out;
  wire par_done_reg1449_done;
  wire par_done_reg1450_in;
  wire par_done_reg1450_write_en;
  wire par_done_reg1450_clk;
  wire par_done_reg1450_out;
  wire par_done_reg1450_done;
  wire par_done_reg1451_in;
  wire par_done_reg1451_write_en;
  wire par_done_reg1451_clk;
  wire par_done_reg1451_out;
  wire par_done_reg1451_done;
  wire par_done_reg1452_in;
  wire par_done_reg1452_write_en;
  wire par_done_reg1452_clk;
  wire par_done_reg1452_out;
  wire par_done_reg1452_done;
  wire par_done_reg1453_in;
  wire par_done_reg1453_write_en;
  wire par_done_reg1453_clk;
  wire par_done_reg1453_out;
  wire par_done_reg1453_done;
  wire par_done_reg1454_in;
  wire par_done_reg1454_write_en;
  wire par_done_reg1454_clk;
  wire par_done_reg1454_out;
  wire par_done_reg1454_done;
  wire par_done_reg1455_in;
  wire par_done_reg1455_write_en;
  wire par_done_reg1455_clk;
  wire par_done_reg1455_out;
  wire par_done_reg1455_done;
  wire par_done_reg1456_in;
  wire par_done_reg1456_write_en;
  wire par_done_reg1456_clk;
  wire par_done_reg1456_out;
  wire par_done_reg1456_done;
  wire par_done_reg1457_in;
  wire par_done_reg1457_write_en;
  wire par_done_reg1457_clk;
  wire par_done_reg1457_out;
  wire par_done_reg1457_done;
  wire par_done_reg1458_in;
  wire par_done_reg1458_write_en;
  wire par_done_reg1458_clk;
  wire par_done_reg1458_out;
  wire par_done_reg1458_done;
  wire par_done_reg1459_in;
  wire par_done_reg1459_write_en;
  wire par_done_reg1459_clk;
  wire par_done_reg1459_out;
  wire par_done_reg1459_done;
  wire par_done_reg1460_in;
  wire par_done_reg1460_write_en;
  wire par_done_reg1460_clk;
  wire par_done_reg1460_out;
  wire par_done_reg1460_done;
  wire par_done_reg1461_in;
  wire par_done_reg1461_write_en;
  wire par_done_reg1461_clk;
  wire par_done_reg1461_out;
  wire par_done_reg1461_done;
  wire par_done_reg1462_in;
  wire par_done_reg1462_write_en;
  wire par_done_reg1462_clk;
  wire par_done_reg1462_out;
  wire par_done_reg1462_done;
  wire par_done_reg1463_in;
  wire par_done_reg1463_write_en;
  wire par_done_reg1463_clk;
  wire par_done_reg1463_out;
  wire par_done_reg1463_done;
  wire par_done_reg1464_in;
  wire par_done_reg1464_write_en;
  wire par_done_reg1464_clk;
  wire par_done_reg1464_out;
  wire par_done_reg1464_done;
  wire par_done_reg1465_in;
  wire par_done_reg1465_write_en;
  wire par_done_reg1465_clk;
  wire par_done_reg1465_out;
  wire par_done_reg1465_done;
  wire par_done_reg1466_in;
  wire par_done_reg1466_write_en;
  wire par_done_reg1466_clk;
  wire par_done_reg1466_out;
  wire par_done_reg1466_done;
  wire par_done_reg1467_in;
  wire par_done_reg1467_write_en;
  wire par_done_reg1467_clk;
  wire par_done_reg1467_out;
  wire par_done_reg1467_done;
  wire par_done_reg1468_in;
  wire par_done_reg1468_write_en;
  wire par_done_reg1468_clk;
  wire par_done_reg1468_out;
  wire par_done_reg1468_done;
  wire par_done_reg1469_in;
  wire par_done_reg1469_write_en;
  wire par_done_reg1469_clk;
  wire par_done_reg1469_out;
  wire par_done_reg1469_done;
  wire par_done_reg1470_in;
  wire par_done_reg1470_write_en;
  wire par_done_reg1470_clk;
  wire par_done_reg1470_out;
  wire par_done_reg1470_done;
  wire par_done_reg1471_in;
  wire par_done_reg1471_write_en;
  wire par_done_reg1471_clk;
  wire par_done_reg1471_out;
  wire par_done_reg1471_done;
  wire par_done_reg1472_in;
  wire par_done_reg1472_write_en;
  wire par_done_reg1472_clk;
  wire par_done_reg1472_out;
  wire par_done_reg1472_done;
  wire par_done_reg1473_in;
  wire par_done_reg1473_write_en;
  wire par_done_reg1473_clk;
  wire par_done_reg1473_out;
  wire par_done_reg1473_done;
  wire par_done_reg1474_in;
  wire par_done_reg1474_write_en;
  wire par_done_reg1474_clk;
  wire par_done_reg1474_out;
  wire par_done_reg1474_done;
  wire par_done_reg1475_in;
  wire par_done_reg1475_write_en;
  wire par_done_reg1475_clk;
  wire par_done_reg1475_out;
  wire par_done_reg1475_done;
  wire par_done_reg1476_in;
  wire par_done_reg1476_write_en;
  wire par_done_reg1476_clk;
  wire par_done_reg1476_out;
  wire par_done_reg1476_done;
  wire par_done_reg1477_in;
  wire par_done_reg1477_write_en;
  wire par_done_reg1477_clk;
  wire par_done_reg1477_out;
  wire par_done_reg1477_done;
  wire par_done_reg1478_in;
  wire par_done_reg1478_write_en;
  wire par_done_reg1478_clk;
  wire par_done_reg1478_out;
  wire par_done_reg1478_done;
  wire par_done_reg1479_in;
  wire par_done_reg1479_write_en;
  wire par_done_reg1479_clk;
  wire par_done_reg1479_out;
  wire par_done_reg1479_done;
  wire par_done_reg1480_in;
  wire par_done_reg1480_write_en;
  wire par_done_reg1480_clk;
  wire par_done_reg1480_out;
  wire par_done_reg1480_done;
  wire par_done_reg1481_in;
  wire par_done_reg1481_write_en;
  wire par_done_reg1481_clk;
  wire par_done_reg1481_out;
  wire par_done_reg1481_done;
  wire par_done_reg1482_in;
  wire par_done_reg1482_write_en;
  wire par_done_reg1482_clk;
  wire par_done_reg1482_out;
  wire par_done_reg1482_done;
  wire par_done_reg1483_in;
  wire par_done_reg1483_write_en;
  wire par_done_reg1483_clk;
  wire par_done_reg1483_out;
  wire par_done_reg1483_done;
  wire par_reset33_in;
  wire par_reset33_write_en;
  wire par_reset33_clk;
  wire par_reset33_out;
  wire par_reset33_done;
  wire par_done_reg1484_in;
  wire par_done_reg1484_write_en;
  wire par_done_reg1484_clk;
  wire par_done_reg1484_out;
  wire par_done_reg1484_done;
  wire par_done_reg1485_in;
  wire par_done_reg1485_write_en;
  wire par_done_reg1485_clk;
  wire par_done_reg1485_out;
  wire par_done_reg1485_done;
  wire par_done_reg1486_in;
  wire par_done_reg1486_write_en;
  wire par_done_reg1486_clk;
  wire par_done_reg1486_out;
  wire par_done_reg1486_done;
  wire par_done_reg1487_in;
  wire par_done_reg1487_write_en;
  wire par_done_reg1487_clk;
  wire par_done_reg1487_out;
  wire par_done_reg1487_done;
  wire par_done_reg1488_in;
  wire par_done_reg1488_write_en;
  wire par_done_reg1488_clk;
  wire par_done_reg1488_out;
  wire par_done_reg1488_done;
  wire par_done_reg1489_in;
  wire par_done_reg1489_write_en;
  wire par_done_reg1489_clk;
  wire par_done_reg1489_out;
  wire par_done_reg1489_done;
  wire par_done_reg1490_in;
  wire par_done_reg1490_write_en;
  wire par_done_reg1490_clk;
  wire par_done_reg1490_out;
  wire par_done_reg1490_done;
  wire par_done_reg1491_in;
  wire par_done_reg1491_write_en;
  wire par_done_reg1491_clk;
  wire par_done_reg1491_out;
  wire par_done_reg1491_done;
  wire par_done_reg1492_in;
  wire par_done_reg1492_write_en;
  wire par_done_reg1492_clk;
  wire par_done_reg1492_out;
  wire par_done_reg1492_done;
  wire par_done_reg1493_in;
  wire par_done_reg1493_write_en;
  wire par_done_reg1493_clk;
  wire par_done_reg1493_out;
  wire par_done_reg1493_done;
  wire par_done_reg1494_in;
  wire par_done_reg1494_write_en;
  wire par_done_reg1494_clk;
  wire par_done_reg1494_out;
  wire par_done_reg1494_done;
  wire par_done_reg1495_in;
  wire par_done_reg1495_write_en;
  wire par_done_reg1495_clk;
  wire par_done_reg1495_out;
  wire par_done_reg1495_done;
  wire par_done_reg1496_in;
  wire par_done_reg1496_write_en;
  wire par_done_reg1496_clk;
  wire par_done_reg1496_out;
  wire par_done_reg1496_done;
  wire par_done_reg1497_in;
  wire par_done_reg1497_write_en;
  wire par_done_reg1497_clk;
  wire par_done_reg1497_out;
  wire par_done_reg1497_done;
  wire par_done_reg1498_in;
  wire par_done_reg1498_write_en;
  wire par_done_reg1498_clk;
  wire par_done_reg1498_out;
  wire par_done_reg1498_done;
  wire par_done_reg1499_in;
  wire par_done_reg1499_write_en;
  wire par_done_reg1499_clk;
  wire par_done_reg1499_out;
  wire par_done_reg1499_done;
  wire par_done_reg1500_in;
  wire par_done_reg1500_write_en;
  wire par_done_reg1500_clk;
  wire par_done_reg1500_out;
  wire par_done_reg1500_done;
  wire par_done_reg1501_in;
  wire par_done_reg1501_write_en;
  wire par_done_reg1501_clk;
  wire par_done_reg1501_out;
  wire par_done_reg1501_done;
  wire par_done_reg1502_in;
  wire par_done_reg1502_write_en;
  wire par_done_reg1502_clk;
  wire par_done_reg1502_out;
  wire par_done_reg1502_done;
  wire par_done_reg1503_in;
  wire par_done_reg1503_write_en;
  wire par_done_reg1503_clk;
  wire par_done_reg1503_out;
  wire par_done_reg1503_done;
  wire par_done_reg1504_in;
  wire par_done_reg1504_write_en;
  wire par_done_reg1504_clk;
  wire par_done_reg1504_out;
  wire par_done_reg1504_done;
  wire par_done_reg1505_in;
  wire par_done_reg1505_write_en;
  wire par_done_reg1505_clk;
  wire par_done_reg1505_out;
  wire par_done_reg1505_done;
  wire par_done_reg1506_in;
  wire par_done_reg1506_write_en;
  wire par_done_reg1506_clk;
  wire par_done_reg1506_out;
  wire par_done_reg1506_done;
  wire par_done_reg1507_in;
  wire par_done_reg1507_write_en;
  wire par_done_reg1507_clk;
  wire par_done_reg1507_out;
  wire par_done_reg1507_done;
  wire par_done_reg1508_in;
  wire par_done_reg1508_write_en;
  wire par_done_reg1508_clk;
  wire par_done_reg1508_out;
  wire par_done_reg1508_done;
  wire par_done_reg1509_in;
  wire par_done_reg1509_write_en;
  wire par_done_reg1509_clk;
  wire par_done_reg1509_out;
  wire par_done_reg1509_done;
  wire par_done_reg1510_in;
  wire par_done_reg1510_write_en;
  wire par_done_reg1510_clk;
  wire par_done_reg1510_out;
  wire par_done_reg1510_done;
  wire par_done_reg1511_in;
  wire par_done_reg1511_write_en;
  wire par_done_reg1511_clk;
  wire par_done_reg1511_out;
  wire par_done_reg1511_done;
  wire par_reset34_in;
  wire par_reset34_write_en;
  wire par_reset34_clk;
  wire par_reset34_out;
  wire par_reset34_done;
  wire par_done_reg1512_in;
  wire par_done_reg1512_write_en;
  wire par_done_reg1512_clk;
  wire par_done_reg1512_out;
  wire par_done_reg1512_done;
  wire par_done_reg1513_in;
  wire par_done_reg1513_write_en;
  wire par_done_reg1513_clk;
  wire par_done_reg1513_out;
  wire par_done_reg1513_done;
  wire par_done_reg1514_in;
  wire par_done_reg1514_write_en;
  wire par_done_reg1514_clk;
  wire par_done_reg1514_out;
  wire par_done_reg1514_done;
  wire par_done_reg1515_in;
  wire par_done_reg1515_write_en;
  wire par_done_reg1515_clk;
  wire par_done_reg1515_out;
  wire par_done_reg1515_done;
  wire par_done_reg1516_in;
  wire par_done_reg1516_write_en;
  wire par_done_reg1516_clk;
  wire par_done_reg1516_out;
  wire par_done_reg1516_done;
  wire par_done_reg1517_in;
  wire par_done_reg1517_write_en;
  wire par_done_reg1517_clk;
  wire par_done_reg1517_out;
  wire par_done_reg1517_done;
  wire par_done_reg1518_in;
  wire par_done_reg1518_write_en;
  wire par_done_reg1518_clk;
  wire par_done_reg1518_out;
  wire par_done_reg1518_done;
  wire par_done_reg1519_in;
  wire par_done_reg1519_write_en;
  wire par_done_reg1519_clk;
  wire par_done_reg1519_out;
  wire par_done_reg1519_done;
  wire par_done_reg1520_in;
  wire par_done_reg1520_write_en;
  wire par_done_reg1520_clk;
  wire par_done_reg1520_out;
  wire par_done_reg1520_done;
  wire par_done_reg1521_in;
  wire par_done_reg1521_write_en;
  wire par_done_reg1521_clk;
  wire par_done_reg1521_out;
  wire par_done_reg1521_done;
  wire par_done_reg1522_in;
  wire par_done_reg1522_write_en;
  wire par_done_reg1522_clk;
  wire par_done_reg1522_out;
  wire par_done_reg1522_done;
  wire par_done_reg1523_in;
  wire par_done_reg1523_write_en;
  wire par_done_reg1523_clk;
  wire par_done_reg1523_out;
  wire par_done_reg1523_done;
  wire par_done_reg1524_in;
  wire par_done_reg1524_write_en;
  wire par_done_reg1524_clk;
  wire par_done_reg1524_out;
  wire par_done_reg1524_done;
  wire par_done_reg1525_in;
  wire par_done_reg1525_write_en;
  wire par_done_reg1525_clk;
  wire par_done_reg1525_out;
  wire par_done_reg1525_done;
  wire par_done_reg1526_in;
  wire par_done_reg1526_write_en;
  wire par_done_reg1526_clk;
  wire par_done_reg1526_out;
  wire par_done_reg1526_done;
  wire par_done_reg1527_in;
  wire par_done_reg1527_write_en;
  wire par_done_reg1527_clk;
  wire par_done_reg1527_out;
  wire par_done_reg1527_done;
  wire par_done_reg1528_in;
  wire par_done_reg1528_write_en;
  wire par_done_reg1528_clk;
  wire par_done_reg1528_out;
  wire par_done_reg1528_done;
  wire par_done_reg1529_in;
  wire par_done_reg1529_write_en;
  wire par_done_reg1529_clk;
  wire par_done_reg1529_out;
  wire par_done_reg1529_done;
  wire par_done_reg1530_in;
  wire par_done_reg1530_write_en;
  wire par_done_reg1530_clk;
  wire par_done_reg1530_out;
  wire par_done_reg1530_done;
  wire par_done_reg1531_in;
  wire par_done_reg1531_write_en;
  wire par_done_reg1531_clk;
  wire par_done_reg1531_out;
  wire par_done_reg1531_done;
  wire par_done_reg1532_in;
  wire par_done_reg1532_write_en;
  wire par_done_reg1532_clk;
  wire par_done_reg1532_out;
  wire par_done_reg1532_done;
  wire par_done_reg1533_in;
  wire par_done_reg1533_write_en;
  wire par_done_reg1533_clk;
  wire par_done_reg1533_out;
  wire par_done_reg1533_done;
  wire par_done_reg1534_in;
  wire par_done_reg1534_write_en;
  wire par_done_reg1534_clk;
  wire par_done_reg1534_out;
  wire par_done_reg1534_done;
  wire par_done_reg1535_in;
  wire par_done_reg1535_write_en;
  wire par_done_reg1535_clk;
  wire par_done_reg1535_out;
  wire par_done_reg1535_done;
  wire par_done_reg1536_in;
  wire par_done_reg1536_write_en;
  wire par_done_reg1536_clk;
  wire par_done_reg1536_out;
  wire par_done_reg1536_done;
  wire par_done_reg1537_in;
  wire par_done_reg1537_write_en;
  wire par_done_reg1537_clk;
  wire par_done_reg1537_out;
  wire par_done_reg1537_done;
  wire par_done_reg1538_in;
  wire par_done_reg1538_write_en;
  wire par_done_reg1538_clk;
  wire par_done_reg1538_out;
  wire par_done_reg1538_done;
  wire par_done_reg1539_in;
  wire par_done_reg1539_write_en;
  wire par_done_reg1539_clk;
  wire par_done_reg1539_out;
  wire par_done_reg1539_done;
  wire par_done_reg1540_in;
  wire par_done_reg1540_write_en;
  wire par_done_reg1540_clk;
  wire par_done_reg1540_out;
  wire par_done_reg1540_done;
  wire par_done_reg1541_in;
  wire par_done_reg1541_write_en;
  wire par_done_reg1541_clk;
  wire par_done_reg1541_out;
  wire par_done_reg1541_done;
  wire par_done_reg1542_in;
  wire par_done_reg1542_write_en;
  wire par_done_reg1542_clk;
  wire par_done_reg1542_out;
  wire par_done_reg1542_done;
  wire par_done_reg1543_in;
  wire par_done_reg1543_write_en;
  wire par_done_reg1543_clk;
  wire par_done_reg1543_out;
  wire par_done_reg1543_done;
  wire par_done_reg1544_in;
  wire par_done_reg1544_write_en;
  wire par_done_reg1544_clk;
  wire par_done_reg1544_out;
  wire par_done_reg1544_done;
  wire par_done_reg1545_in;
  wire par_done_reg1545_write_en;
  wire par_done_reg1545_clk;
  wire par_done_reg1545_out;
  wire par_done_reg1545_done;
  wire par_done_reg1546_in;
  wire par_done_reg1546_write_en;
  wire par_done_reg1546_clk;
  wire par_done_reg1546_out;
  wire par_done_reg1546_done;
  wire par_done_reg1547_in;
  wire par_done_reg1547_write_en;
  wire par_done_reg1547_clk;
  wire par_done_reg1547_out;
  wire par_done_reg1547_done;
  wire par_done_reg1548_in;
  wire par_done_reg1548_write_en;
  wire par_done_reg1548_clk;
  wire par_done_reg1548_out;
  wire par_done_reg1548_done;
  wire par_done_reg1549_in;
  wire par_done_reg1549_write_en;
  wire par_done_reg1549_clk;
  wire par_done_reg1549_out;
  wire par_done_reg1549_done;
  wire par_done_reg1550_in;
  wire par_done_reg1550_write_en;
  wire par_done_reg1550_clk;
  wire par_done_reg1550_out;
  wire par_done_reg1550_done;
  wire par_done_reg1551_in;
  wire par_done_reg1551_write_en;
  wire par_done_reg1551_clk;
  wire par_done_reg1551_out;
  wire par_done_reg1551_done;
  wire par_done_reg1552_in;
  wire par_done_reg1552_write_en;
  wire par_done_reg1552_clk;
  wire par_done_reg1552_out;
  wire par_done_reg1552_done;
  wire par_done_reg1553_in;
  wire par_done_reg1553_write_en;
  wire par_done_reg1553_clk;
  wire par_done_reg1553_out;
  wire par_done_reg1553_done;
  wire par_reset35_in;
  wire par_reset35_write_en;
  wire par_reset35_clk;
  wire par_reset35_out;
  wire par_reset35_done;
  wire par_done_reg1554_in;
  wire par_done_reg1554_write_en;
  wire par_done_reg1554_clk;
  wire par_done_reg1554_out;
  wire par_done_reg1554_done;
  wire par_done_reg1555_in;
  wire par_done_reg1555_write_en;
  wire par_done_reg1555_clk;
  wire par_done_reg1555_out;
  wire par_done_reg1555_done;
  wire par_done_reg1556_in;
  wire par_done_reg1556_write_en;
  wire par_done_reg1556_clk;
  wire par_done_reg1556_out;
  wire par_done_reg1556_done;
  wire par_done_reg1557_in;
  wire par_done_reg1557_write_en;
  wire par_done_reg1557_clk;
  wire par_done_reg1557_out;
  wire par_done_reg1557_done;
  wire par_done_reg1558_in;
  wire par_done_reg1558_write_en;
  wire par_done_reg1558_clk;
  wire par_done_reg1558_out;
  wire par_done_reg1558_done;
  wire par_done_reg1559_in;
  wire par_done_reg1559_write_en;
  wire par_done_reg1559_clk;
  wire par_done_reg1559_out;
  wire par_done_reg1559_done;
  wire par_done_reg1560_in;
  wire par_done_reg1560_write_en;
  wire par_done_reg1560_clk;
  wire par_done_reg1560_out;
  wire par_done_reg1560_done;
  wire par_done_reg1561_in;
  wire par_done_reg1561_write_en;
  wire par_done_reg1561_clk;
  wire par_done_reg1561_out;
  wire par_done_reg1561_done;
  wire par_done_reg1562_in;
  wire par_done_reg1562_write_en;
  wire par_done_reg1562_clk;
  wire par_done_reg1562_out;
  wire par_done_reg1562_done;
  wire par_done_reg1563_in;
  wire par_done_reg1563_write_en;
  wire par_done_reg1563_clk;
  wire par_done_reg1563_out;
  wire par_done_reg1563_done;
  wire par_done_reg1564_in;
  wire par_done_reg1564_write_en;
  wire par_done_reg1564_clk;
  wire par_done_reg1564_out;
  wire par_done_reg1564_done;
  wire par_done_reg1565_in;
  wire par_done_reg1565_write_en;
  wire par_done_reg1565_clk;
  wire par_done_reg1565_out;
  wire par_done_reg1565_done;
  wire par_done_reg1566_in;
  wire par_done_reg1566_write_en;
  wire par_done_reg1566_clk;
  wire par_done_reg1566_out;
  wire par_done_reg1566_done;
  wire par_done_reg1567_in;
  wire par_done_reg1567_write_en;
  wire par_done_reg1567_clk;
  wire par_done_reg1567_out;
  wire par_done_reg1567_done;
  wire par_done_reg1568_in;
  wire par_done_reg1568_write_en;
  wire par_done_reg1568_clk;
  wire par_done_reg1568_out;
  wire par_done_reg1568_done;
  wire par_done_reg1569_in;
  wire par_done_reg1569_write_en;
  wire par_done_reg1569_clk;
  wire par_done_reg1569_out;
  wire par_done_reg1569_done;
  wire par_done_reg1570_in;
  wire par_done_reg1570_write_en;
  wire par_done_reg1570_clk;
  wire par_done_reg1570_out;
  wire par_done_reg1570_done;
  wire par_done_reg1571_in;
  wire par_done_reg1571_write_en;
  wire par_done_reg1571_clk;
  wire par_done_reg1571_out;
  wire par_done_reg1571_done;
  wire par_done_reg1572_in;
  wire par_done_reg1572_write_en;
  wire par_done_reg1572_clk;
  wire par_done_reg1572_out;
  wire par_done_reg1572_done;
  wire par_done_reg1573_in;
  wire par_done_reg1573_write_en;
  wire par_done_reg1573_clk;
  wire par_done_reg1573_out;
  wire par_done_reg1573_done;
  wire par_done_reg1574_in;
  wire par_done_reg1574_write_en;
  wire par_done_reg1574_clk;
  wire par_done_reg1574_out;
  wire par_done_reg1574_done;
  wire par_reset36_in;
  wire par_reset36_write_en;
  wire par_reset36_clk;
  wire par_reset36_out;
  wire par_reset36_done;
  wire par_done_reg1575_in;
  wire par_done_reg1575_write_en;
  wire par_done_reg1575_clk;
  wire par_done_reg1575_out;
  wire par_done_reg1575_done;
  wire par_done_reg1576_in;
  wire par_done_reg1576_write_en;
  wire par_done_reg1576_clk;
  wire par_done_reg1576_out;
  wire par_done_reg1576_done;
  wire par_done_reg1577_in;
  wire par_done_reg1577_write_en;
  wire par_done_reg1577_clk;
  wire par_done_reg1577_out;
  wire par_done_reg1577_done;
  wire par_done_reg1578_in;
  wire par_done_reg1578_write_en;
  wire par_done_reg1578_clk;
  wire par_done_reg1578_out;
  wire par_done_reg1578_done;
  wire par_done_reg1579_in;
  wire par_done_reg1579_write_en;
  wire par_done_reg1579_clk;
  wire par_done_reg1579_out;
  wire par_done_reg1579_done;
  wire par_done_reg1580_in;
  wire par_done_reg1580_write_en;
  wire par_done_reg1580_clk;
  wire par_done_reg1580_out;
  wire par_done_reg1580_done;
  wire par_done_reg1581_in;
  wire par_done_reg1581_write_en;
  wire par_done_reg1581_clk;
  wire par_done_reg1581_out;
  wire par_done_reg1581_done;
  wire par_done_reg1582_in;
  wire par_done_reg1582_write_en;
  wire par_done_reg1582_clk;
  wire par_done_reg1582_out;
  wire par_done_reg1582_done;
  wire par_done_reg1583_in;
  wire par_done_reg1583_write_en;
  wire par_done_reg1583_clk;
  wire par_done_reg1583_out;
  wire par_done_reg1583_done;
  wire par_done_reg1584_in;
  wire par_done_reg1584_write_en;
  wire par_done_reg1584_clk;
  wire par_done_reg1584_out;
  wire par_done_reg1584_done;
  wire par_done_reg1585_in;
  wire par_done_reg1585_write_en;
  wire par_done_reg1585_clk;
  wire par_done_reg1585_out;
  wire par_done_reg1585_done;
  wire par_done_reg1586_in;
  wire par_done_reg1586_write_en;
  wire par_done_reg1586_clk;
  wire par_done_reg1586_out;
  wire par_done_reg1586_done;
  wire par_done_reg1587_in;
  wire par_done_reg1587_write_en;
  wire par_done_reg1587_clk;
  wire par_done_reg1587_out;
  wire par_done_reg1587_done;
  wire par_done_reg1588_in;
  wire par_done_reg1588_write_en;
  wire par_done_reg1588_clk;
  wire par_done_reg1588_out;
  wire par_done_reg1588_done;
  wire par_done_reg1589_in;
  wire par_done_reg1589_write_en;
  wire par_done_reg1589_clk;
  wire par_done_reg1589_out;
  wire par_done_reg1589_done;
  wire par_done_reg1590_in;
  wire par_done_reg1590_write_en;
  wire par_done_reg1590_clk;
  wire par_done_reg1590_out;
  wire par_done_reg1590_done;
  wire par_done_reg1591_in;
  wire par_done_reg1591_write_en;
  wire par_done_reg1591_clk;
  wire par_done_reg1591_out;
  wire par_done_reg1591_done;
  wire par_done_reg1592_in;
  wire par_done_reg1592_write_en;
  wire par_done_reg1592_clk;
  wire par_done_reg1592_out;
  wire par_done_reg1592_done;
  wire par_done_reg1593_in;
  wire par_done_reg1593_write_en;
  wire par_done_reg1593_clk;
  wire par_done_reg1593_out;
  wire par_done_reg1593_done;
  wire par_done_reg1594_in;
  wire par_done_reg1594_write_en;
  wire par_done_reg1594_clk;
  wire par_done_reg1594_out;
  wire par_done_reg1594_done;
  wire par_done_reg1595_in;
  wire par_done_reg1595_write_en;
  wire par_done_reg1595_clk;
  wire par_done_reg1595_out;
  wire par_done_reg1595_done;
  wire par_done_reg1596_in;
  wire par_done_reg1596_write_en;
  wire par_done_reg1596_clk;
  wire par_done_reg1596_out;
  wire par_done_reg1596_done;
  wire par_done_reg1597_in;
  wire par_done_reg1597_write_en;
  wire par_done_reg1597_clk;
  wire par_done_reg1597_out;
  wire par_done_reg1597_done;
  wire par_done_reg1598_in;
  wire par_done_reg1598_write_en;
  wire par_done_reg1598_clk;
  wire par_done_reg1598_out;
  wire par_done_reg1598_done;
  wire par_done_reg1599_in;
  wire par_done_reg1599_write_en;
  wire par_done_reg1599_clk;
  wire par_done_reg1599_out;
  wire par_done_reg1599_done;
  wire par_done_reg1600_in;
  wire par_done_reg1600_write_en;
  wire par_done_reg1600_clk;
  wire par_done_reg1600_out;
  wire par_done_reg1600_done;
  wire par_done_reg1601_in;
  wire par_done_reg1601_write_en;
  wire par_done_reg1601_clk;
  wire par_done_reg1601_out;
  wire par_done_reg1601_done;
  wire par_done_reg1602_in;
  wire par_done_reg1602_write_en;
  wire par_done_reg1602_clk;
  wire par_done_reg1602_out;
  wire par_done_reg1602_done;
  wire par_done_reg1603_in;
  wire par_done_reg1603_write_en;
  wire par_done_reg1603_clk;
  wire par_done_reg1603_out;
  wire par_done_reg1603_done;
  wire par_done_reg1604_in;
  wire par_done_reg1604_write_en;
  wire par_done_reg1604_clk;
  wire par_done_reg1604_out;
  wire par_done_reg1604_done;
  wire par_reset37_in;
  wire par_reset37_write_en;
  wire par_reset37_clk;
  wire par_reset37_out;
  wire par_reset37_done;
  wire par_done_reg1605_in;
  wire par_done_reg1605_write_en;
  wire par_done_reg1605_clk;
  wire par_done_reg1605_out;
  wire par_done_reg1605_done;
  wire par_done_reg1606_in;
  wire par_done_reg1606_write_en;
  wire par_done_reg1606_clk;
  wire par_done_reg1606_out;
  wire par_done_reg1606_done;
  wire par_done_reg1607_in;
  wire par_done_reg1607_write_en;
  wire par_done_reg1607_clk;
  wire par_done_reg1607_out;
  wire par_done_reg1607_done;
  wire par_done_reg1608_in;
  wire par_done_reg1608_write_en;
  wire par_done_reg1608_clk;
  wire par_done_reg1608_out;
  wire par_done_reg1608_done;
  wire par_done_reg1609_in;
  wire par_done_reg1609_write_en;
  wire par_done_reg1609_clk;
  wire par_done_reg1609_out;
  wire par_done_reg1609_done;
  wire par_done_reg1610_in;
  wire par_done_reg1610_write_en;
  wire par_done_reg1610_clk;
  wire par_done_reg1610_out;
  wire par_done_reg1610_done;
  wire par_done_reg1611_in;
  wire par_done_reg1611_write_en;
  wire par_done_reg1611_clk;
  wire par_done_reg1611_out;
  wire par_done_reg1611_done;
  wire par_done_reg1612_in;
  wire par_done_reg1612_write_en;
  wire par_done_reg1612_clk;
  wire par_done_reg1612_out;
  wire par_done_reg1612_done;
  wire par_done_reg1613_in;
  wire par_done_reg1613_write_en;
  wire par_done_reg1613_clk;
  wire par_done_reg1613_out;
  wire par_done_reg1613_done;
  wire par_done_reg1614_in;
  wire par_done_reg1614_write_en;
  wire par_done_reg1614_clk;
  wire par_done_reg1614_out;
  wire par_done_reg1614_done;
  wire par_done_reg1615_in;
  wire par_done_reg1615_write_en;
  wire par_done_reg1615_clk;
  wire par_done_reg1615_out;
  wire par_done_reg1615_done;
  wire par_done_reg1616_in;
  wire par_done_reg1616_write_en;
  wire par_done_reg1616_clk;
  wire par_done_reg1616_out;
  wire par_done_reg1616_done;
  wire par_done_reg1617_in;
  wire par_done_reg1617_write_en;
  wire par_done_reg1617_clk;
  wire par_done_reg1617_out;
  wire par_done_reg1617_done;
  wire par_done_reg1618_in;
  wire par_done_reg1618_write_en;
  wire par_done_reg1618_clk;
  wire par_done_reg1618_out;
  wire par_done_reg1618_done;
  wire par_done_reg1619_in;
  wire par_done_reg1619_write_en;
  wire par_done_reg1619_clk;
  wire par_done_reg1619_out;
  wire par_done_reg1619_done;
  wire par_reset38_in;
  wire par_reset38_write_en;
  wire par_reset38_clk;
  wire par_reset38_out;
  wire par_reset38_done;
  wire par_done_reg1620_in;
  wire par_done_reg1620_write_en;
  wire par_done_reg1620_clk;
  wire par_done_reg1620_out;
  wire par_done_reg1620_done;
  wire par_done_reg1621_in;
  wire par_done_reg1621_write_en;
  wire par_done_reg1621_clk;
  wire par_done_reg1621_out;
  wire par_done_reg1621_done;
  wire par_done_reg1622_in;
  wire par_done_reg1622_write_en;
  wire par_done_reg1622_clk;
  wire par_done_reg1622_out;
  wire par_done_reg1622_done;
  wire par_done_reg1623_in;
  wire par_done_reg1623_write_en;
  wire par_done_reg1623_clk;
  wire par_done_reg1623_out;
  wire par_done_reg1623_done;
  wire par_done_reg1624_in;
  wire par_done_reg1624_write_en;
  wire par_done_reg1624_clk;
  wire par_done_reg1624_out;
  wire par_done_reg1624_done;
  wire par_done_reg1625_in;
  wire par_done_reg1625_write_en;
  wire par_done_reg1625_clk;
  wire par_done_reg1625_out;
  wire par_done_reg1625_done;
  wire par_done_reg1626_in;
  wire par_done_reg1626_write_en;
  wire par_done_reg1626_clk;
  wire par_done_reg1626_out;
  wire par_done_reg1626_done;
  wire par_done_reg1627_in;
  wire par_done_reg1627_write_en;
  wire par_done_reg1627_clk;
  wire par_done_reg1627_out;
  wire par_done_reg1627_done;
  wire par_done_reg1628_in;
  wire par_done_reg1628_write_en;
  wire par_done_reg1628_clk;
  wire par_done_reg1628_out;
  wire par_done_reg1628_done;
  wire par_done_reg1629_in;
  wire par_done_reg1629_write_en;
  wire par_done_reg1629_clk;
  wire par_done_reg1629_out;
  wire par_done_reg1629_done;
  wire par_done_reg1630_in;
  wire par_done_reg1630_write_en;
  wire par_done_reg1630_clk;
  wire par_done_reg1630_out;
  wire par_done_reg1630_done;
  wire par_done_reg1631_in;
  wire par_done_reg1631_write_en;
  wire par_done_reg1631_clk;
  wire par_done_reg1631_out;
  wire par_done_reg1631_done;
  wire par_done_reg1632_in;
  wire par_done_reg1632_write_en;
  wire par_done_reg1632_clk;
  wire par_done_reg1632_out;
  wire par_done_reg1632_done;
  wire par_done_reg1633_in;
  wire par_done_reg1633_write_en;
  wire par_done_reg1633_clk;
  wire par_done_reg1633_out;
  wire par_done_reg1633_done;
  wire par_done_reg1634_in;
  wire par_done_reg1634_write_en;
  wire par_done_reg1634_clk;
  wire par_done_reg1634_out;
  wire par_done_reg1634_done;
  wire par_done_reg1635_in;
  wire par_done_reg1635_write_en;
  wire par_done_reg1635_clk;
  wire par_done_reg1635_out;
  wire par_done_reg1635_done;
  wire par_done_reg1636_in;
  wire par_done_reg1636_write_en;
  wire par_done_reg1636_clk;
  wire par_done_reg1636_out;
  wire par_done_reg1636_done;
  wire par_done_reg1637_in;
  wire par_done_reg1637_write_en;
  wire par_done_reg1637_clk;
  wire par_done_reg1637_out;
  wire par_done_reg1637_done;
  wire par_done_reg1638_in;
  wire par_done_reg1638_write_en;
  wire par_done_reg1638_clk;
  wire par_done_reg1638_out;
  wire par_done_reg1638_done;
  wire par_done_reg1639_in;
  wire par_done_reg1639_write_en;
  wire par_done_reg1639_clk;
  wire par_done_reg1639_out;
  wire par_done_reg1639_done;
  wire par_reset39_in;
  wire par_reset39_write_en;
  wire par_reset39_clk;
  wire par_reset39_out;
  wire par_reset39_done;
  wire par_done_reg1640_in;
  wire par_done_reg1640_write_en;
  wire par_done_reg1640_clk;
  wire par_done_reg1640_out;
  wire par_done_reg1640_done;
  wire par_done_reg1641_in;
  wire par_done_reg1641_write_en;
  wire par_done_reg1641_clk;
  wire par_done_reg1641_out;
  wire par_done_reg1641_done;
  wire par_done_reg1642_in;
  wire par_done_reg1642_write_en;
  wire par_done_reg1642_clk;
  wire par_done_reg1642_out;
  wire par_done_reg1642_done;
  wire par_done_reg1643_in;
  wire par_done_reg1643_write_en;
  wire par_done_reg1643_clk;
  wire par_done_reg1643_out;
  wire par_done_reg1643_done;
  wire par_done_reg1644_in;
  wire par_done_reg1644_write_en;
  wire par_done_reg1644_clk;
  wire par_done_reg1644_out;
  wire par_done_reg1644_done;
  wire par_done_reg1645_in;
  wire par_done_reg1645_write_en;
  wire par_done_reg1645_clk;
  wire par_done_reg1645_out;
  wire par_done_reg1645_done;
  wire par_done_reg1646_in;
  wire par_done_reg1646_write_en;
  wire par_done_reg1646_clk;
  wire par_done_reg1646_out;
  wire par_done_reg1646_done;
  wire par_done_reg1647_in;
  wire par_done_reg1647_write_en;
  wire par_done_reg1647_clk;
  wire par_done_reg1647_out;
  wire par_done_reg1647_done;
  wire par_done_reg1648_in;
  wire par_done_reg1648_write_en;
  wire par_done_reg1648_clk;
  wire par_done_reg1648_out;
  wire par_done_reg1648_done;
  wire par_done_reg1649_in;
  wire par_done_reg1649_write_en;
  wire par_done_reg1649_clk;
  wire par_done_reg1649_out;
  wire par_done_reg1649_done;
  wire par_reset40_in;
  wire par_reset40_write_en;
  wire par_reset40_clk;
  wire par_reset40_out;
  wire par_reset40_done;
  wire par_done_reg1650_in;
  wire par_done_reg1650_write_en;
  wire par_done_reg1650_clk;
  wire par_done_reg1650_out;
  wire par_done_reg1650_done;
  wire par_done_reg1651_in;
  wire par_done_reg1651_write_en;
  wire par_done_reg1651_clk;
  wire par_done_reg1651_out;
  wire par_done_reg1651_done;
  wire par_done_reg1652_in;
  wire par_done_reg1652_write_en;
  wire par_done_reg1652_clk;
  wire par_done_reg1652_out;
  wire par_done_reg1652_done;
  wire par_done_reg1653_in;
  wire par_done_reg1653_write_en;
  wire par_done_reg1653_clk;
  wire par_done_reg1653_out;
  wire par_done_reg1653_done;
  wire par_done_reg1654_in;
  wire par_done_reg1654_write_en;
  wire par_done_reg1654_clk;
  wire par_done_reg1654_out;
  wire par_done_reg1654_done;
  wire par_done_reg1655_in;
  wire par_done_reg1655_write_en;
  wire par_done_reg1655_clk;
  wire par_done_reg1655_out;
  wire par_done_reg1655_done;
  wire par_done_reg1656_in;
  wire par_done_reg1656_write_en;
  wire par_done_reg1656_clk;
  wire par_done_reg1656_out;
  wire par_done_reg1656_done;
  wire par_done_reg1657_in;
  wire par_done_reg1657_write_en;
  wire par_done_reg1657_clk;
  wire par_done_reg1657_out;
  wire par_done_reg1657_done;
  wire par_done_reg1658_in;
  wire par_done_reg1658_write_en;
  wire par_done_reg1658_clk;
  wire par_done_reg1658_out;
  wire par_done_reg1658_done;
  wire par_done_reg1659_in;
  wire par_done_reg1659_write_en;
  wire par_done_reg1659_clk;
  wire par_done_reg1659_out;
  wire par_done_reg1659_done;
  wire par_done_reg1660_in;
  wire par_done_reg1660_write_en;
  wire par_done_reg1660_clk;
  wire par_done_reg1660_out;
  wire par_done_reg1660_done;
  wire par_done_reg1661_in;
  wire par_done_reg1661_write_en;
  wire par_done_reg1661_clk;
  wire par_done_reg1661_out;
  wire par_done_reg1661_done;
  wire par_reset41_in;
  wire par_reset41_write_en;
  wire par_reset41_clk;
  wire par_reset41_out;
  wire par_reset41_done;
  wire par_done_reg1662_in;
  wire par_done_reg1662_write_en;
  wire par_done_reg1662_clk;
  wire par_done_reg1662_out;
  wire par_done_reg1662_done;
  wire par_done_reg1663_in;
  wire par_done_reg1663_write_en;
  wire par_done_reg1663_clk;
  wire par_done_reg1663_out;
  wire par_done_reg1663_done;
  wire par_done_reg1664_in;
  wire par_done_reg1664_write_en;
  wire par_done_reg1664_clk;
  wire par_done_reg1664_out;
  wire par_done_reg1664_done;
  wire par_done_reg1665_in;
  wire par_done_reg1665_write_en;
  wire par_done_reg1665_clk;
  wire par_done_reg1665_out;
  wire par_done_reg1665_done;
  wire par_done_reg1666_in;
  wire par_done_reg1666_write_en;
  wire par_done_reg1666_clk;
  wire par_done_reg1666_out;
  wire par_done_reg1666_done;
  wire par_done_reg1667_in;
  wire par_done_reg1667_write_en;
  wire par_done_reg1667_clk;
  wire par_done_reg1667_out;
  wire par_done_reg1667_done;
  wire par_reset42_in;
  wire par_reset42_write_en;
  wire par_reset42_clk;
  wire par_reset42_out;
  wire par_reset42_done;
  wire par_done_reg1668_in;
  wire par_done_reg1668_write_en;
  wire par_done_reg1668_clk;
  wire par_done_reg1668_out;
  wire par_done_reg1668_done;
  wire par_done_reg1669_in;
  wire par_done_reg1669_write_en;
  wire par_done_reg1669_clk;
  wire par_done_reg1669_out;
  wire par_done_reg1669_done;
  wire par_done_reg1670_in;
  wire par_done_reg1670_write_en;
  wire par_done_reg1670_clk;
  wire par_done_reg1670_out;
  wire par_done_reg1670_done;
  wire par_done_reg1671_in;
  wire par_done_reg1671_write_en;
  wire par_done_reg1671_clk;
  wire par_done_reg1671_out;
  wire par_done_reg1671_done;
  wire par_done_reg1672_in;
  wire par_done_reg1672_write_en;
  wire par_done_reg1672_clk;
  wire par_done_reg1672_out;
  wire par_done_reg1672_done;
  wire par_done_reg1673_in;
  wire par_done_reg1673_write_en;
  wire par_done_reg1673_clk;
  wire par_done_reg1673_out;
  wire par_done_reg1673_done;
  wire par_reset43_in;
  wire par_reset43_write_en;
  wire par_reset43_clk;
  wire par_reset43_out;
  wire par_reset43_done;
  wire par_done_reg1674_in;
  wire par_done_reg1674_write_en;
  wire par_done_reg1674_clk;
  wire par_done_reg1674_out;
  wire par_done_reg1674_done;
  wire par_done_reg1675_in;
  wire par_done_reg1675_write_en;
  wire par_done_reg1675_clk;
  wire par_done_reg1675_out;
  wire par_done_reg1675_done;
  wire par_done_reg1676_in;
  wire par_done_reg1676_write_en;
  wire par_done_reg1676_clk;
  wire par_done_reg1676_out;
  wire par_done_reg1676_done;
  wire par_reset44_in;
  wire par_reset44_write_en;
  wire par_reset44_clk;
  wire par_reset44_out;
  wire par_reset44_done;
  wire par_done_reg1677_in;
  wire par_done_reg1677_write_en;
  wire par_done_reg1677_clk;
  wire par_done_reg1677_out;
  wire par_done_reg1677_done;
  wire par_done_reg1678_in;
  wire par_done_reg1678_write_en;
  wire par_done_reg1678_clk;
  wire par_done_reg1678_out;
  wire par_done_reg1678_done;
  wire par_reset45_in;
  wire par_reset45_write_en;
  wire par_reset45_clk;
  wire par_reset45_out;
  wire par_reset45_done;
  wire par_done_reg1679_in;
  wire par_done_reg1679_write_en;
  wire par_done_reg1679_clk;
  wire par_done_reg1679_out;
  wire par_done_reg1679_done;
  wire [31:0] fsm0_in;
  wire fsm0_write_en;
  wire fsm0_clk;
  wire [31:0] fsm0_out;
  wire fsm0_done;
  
  // Subcomponent Instances
  std_reg #(32) left_77_read (
      .in(left_77_read_in),
      .write_en(left_77_read_write_en),
      .clk(clk),
      .out(left_77_read_out),
      .done(left_77_read_done)
  );
  
  std_reg #(32) top_77_read (
      .in(top_77_read_in),
      .write_en(top_77_read_write_en),
      .clk(clk),
      .out(top_77_read_out),
      .done(top_77_read_done)
  );
  
  mac_pe #() pe_77 (
      .top(pe_77_top),
      .left(pe_77_left),
      .go(pe_77_go),
      .clk(clk),
      .down(pe_77_down),
      .right(pe_77_right),
      .out(pe_77_out),
      .done(pe_77_done)
  );
  
  std_reg #(32) right_76_write (
      .in(right_76_write_in),
      .write_en(right_76_write_write_en),
      .clk(clk),
      .out(right_76_write_out),
      .done(right_76_write_done)
  );
  
  std_reg #(32) left_76_read (
      .in(left_76_read_in),
      .write_en(left_76_read_write_en),
      .clk(clk),
      .out(left_76_read_out),
      .done(left_76_read_done)
  );
  
  std_reg #(32) top_76_read (
      .in(top_76_read_in),
      .write_en(top_76_read_write_en),
      .clk(clk),
      .out(top_76_read_out),
      .done(top_76_read_done)
  );
  
  mac_pe #() pe_76 (
      .top(pe_76_top),
      .left(pe_76_left),
      .go(pe_76_go),
      .clk(clk),
      .down(pe_76_down),
      .right(pe_76_right),
      .out(pe_76_out),
      .done(pe_76_done)
  );
  
  std_reg #(32) right_75_write (
      .in(right_75_write_in),
      .write_en(right_75_write_write_en),
      .clk(clk),
      .out(right_75_write_out),
      .done(right_75_write_done)
  );
  
  std_reg #(32) left_75_read (
      .in(left_75_read_in),
      .write_en(left_75_read_write_en),
      .clk(clk),
      .out(left_75_read_out),
      .done(left_75_read_done)
  );
  
  std_reg #(32) top_75_read (
      .in(top_75_read_in),
      .write_en(top_75_read_write_en),
      .clk(clk),
      .out(top_75_read_out),
      .done(top_75_read_done)
  );
  
  mac_pe #() pe_75 (
      .top(pe_75_top),
      .left(pe_75_left),
      .go(pe_75_go),
      .clk(clk),
      .down(pe_75_down),
      .right(pe_75_right),
      .out(pe_75_out),
      .done(pe_75_done)
  );
  
  std_reg #(32) right_74_write (
      .in(right_74_write_in),
      .write_en(right_74_write_write_en),
      .clk(clk),
      .out(right_74_write_out),
      .done(right_74_write_done)
  );
  
  std_reg #(32) left_74_read (
      .in(left_74_read_in),
      .write_en(left_74_read_write_en),
      .clk(clk),
      .out(left_74_read_out),
      .done(left_74_read_done)
  );
  
  std_reg #(32) top_74_read (
      .in(top_74_read_in),
      .write_en(top_74_read_write_en),
      .clk(clk),
      .out(top_74_read_out),
      .done(top_74_read_done)
  );
  
  mac_pe #() pe_74 (
      .top(pe_74_top),
      .left(pe_74_left),
      .go(pe_74_go),
      .clk(clk),
      .down(pe_74_down),
      .right(pe_74_right),
      .out(pe_74_out),
      .done(pe_74_done)
  );
  
  std_reg #(32) right_73_write (
      .in(right_73_write_in),
      .write_en(right_73_write_write_en),
      .clk(clk),
      .out(right_73_write_out),
      .done(right_73_write_done)
  );
  
  std_reg #(32) left_73_read (
      .in(left_73_read_in),
      .write_en(left_73_read_write_en),
      .clk(clk),
      .out(left_73_read_out),
      .done(left_73_read_done)
  );
  
  std_reg #(32) top_73_read (
      .in(top_73_read_in),
      .write_en(top_73_read_write_en),
      .clk(clk),
      .out(top_73_read_out),
      .done(top_73_read_done)
  );
  
  mac_pe #() pe_73 (
      .top(pe_73_top),
      .left(pe_73_left),
      .go(pe_73_go),
      .clk(clk),
      .down(pe_73_down),
      .right(pe_73_right),
      .out(pe_73_out),
      .done(pe_73_done)
  );
  
  std_reg #(32) right_72_write (
      .in(right_72_write_in),
      .write_en(right_72_write_write_en),
      .clk(clk),
      .out(right_72_write_out),
      .done(right_72_write_done)
  );
  
  std_reg #(32) left_72_read (
      .in(left_72_read_in),
      .write_en(left_72_read_write_en),
      .clk(clk),
      .out(left_72_read_out),
      .done(left_72_read_done)
  );
  
  std_reg #(32) top_72_read (
      .in(top_72_read_in),
      .write_en(top_72_read_write_en),
      .clk(clk),
      .out(top_72_read_out),
      .done(top_72_read_done)
  );
  
  mac_pe #() pe_72 (
      .top(pe_72_top),
      .left(pe_72_left),
      .go(pe_72_go),
      .clk(clk),
      .down(pe_72_down),
      .right(pe_72_right),
      .out(pe_72_out),
      .done(pe_72_done)
  );
  
  std_reg #(32) right_71_write (
      .in(right_71_write_in),
      .write_en(right_71_write_write_en),
      .clk(clk),
      .out(right_71_write_out),
      .done(right_71_write_done)
  );
  
  std_reg #(32) left_71_read (
      .in(left_71_read_in),
      .write_en(left_71_read_write_en),
      .clk(clk),
      .out(left_71_read_out),
      .done(left_71_read_done)
  );
  
  std_reg #(32) top_71_read (
      .in(top_71_read_in),
      .write_en(top_71_read_write_en),
      .clk(clk),
      .out(top_71_read_out),
      .done(top_71_read_done)
  );
  
  mac_pe #() pe_71 (
      .top(pe_71_top),
      .left(pe_71_left),
      .go(pe_71_go),
      .clk(clk),
      .down(pe_71_down),
      .right(pe_71_right),
      .out(pe_71_out),
      .done(pe_71_done)
  );
  
  std_reg #(32) right_70_write (
      .in(right_70_write_in),
      .write_en(right_70_write_write_en),
      .clk(clk),
      .out(right_70_write_out),
      .done(right_70_write_done)
  );
  
  std_reg #(32) left_70_read (
      .in(left_70_read_in),
      .write_en(left_70_read_write_en),
      .clk(clk),
      .out(left_70_read_out),
      .done(left_70_read_done)
  );
  
  std_reg #(32) top_70_read (
      .in(top_70_read_in),
      .write_en(top_70_read_write_en),
      .clk(clk),
      .out(top_70_read_out),
      .done(top_70_read_done)
  );
  
  mac_pe #() pe_70 (
      .top(pe_70_top),
      .left(pe_70_left),
      .go(pe_70_go),
      .clk(clk),
      .down(pe_70_down),
      .right(pe_70_right),
      .out(pe_70_out),
      .done(pe_70_done)
  );
  
  std_reg #(32) down_67_write (
      .in(down_67_write_in),
      .write_en(down_67_write_write_en),
      .clk(clk),
      .out(down_67_write_out),
      .done(down_67_write_done)
  );
  
  std_reg #(32) left_67_read (
      .in(left_67_read_in),
      .write_en(left_67_read_write_en),
      .clk(clk),
      .out(left_67_read_out),
      .done(left_67_read_done)
  );
  
  std_reg #(32) top_67_read (
      .in(top_67_read_in),
      .write_en(top_67_read_write_en),
      .clk(clk),
      .out(top_67_read_out),
      .done(top_67_read_done)
  );
  
  mac_pe #() pe_67 (
      .top(pe_67_top),
      .left(pe_67_left),
      .go(pe_67_go),
      .clk(clk),
      .down(pe_67_down),
      .right(pe_67_right),
      .out(pe_67_out),
      .done(pe_67_done)
  );
  
  std_reg #(32) down_66_write (
      .in(down_66_write_in),
      .write_en(down_66_write_write_en),
      .clk(clk),
      .out(down_66_write_out),
      .done(down_66_write_done)
  );
  
  std_reg #(32) right_66_write (
      .in(right_66_write_in),
      .write_en(right_66_write_write_en),
      .clk(clk),
      .out(right_66_write_out),
      .done(right_66_write_done)
  );
  
  std_reg #(32) left_66_read (
      .in(left_66_read_in),
      .write_en(left_66_read_write_en),
      .clk(clk),
      .out(left_66_read_out),
      .done(left_66_read_done)
  );
  
  std_reg #(32) top_66_read (
      .in(top_66_read_in),
      .write_en(top_66_read_write_en),
      .clk(clk),
      .out(top_66_read_out),
      .done(top_66_read_done)
  );
  
  mac_pe #() pe_66 (
      .top(pe_66_top),
      .left(pe_66_left),
      .go(pe_66_go),
      .clk(clk),
      .down(pe_66_down),
      .right(pe_66_right),
      .out(pe_66_out),
      .done(pe_66_done)
  );
  
  std_reg #(32) down_65_write (
      .in(down_65_write_in),
      .write_en(down_65_write_write_en),
      .clk(clk),
      .out(down_65_write_out),
      .done(down_65_write_done)
  );
  
  std_reg #(32) right_65_write (
      .in(right_65_write_in),
      .write_en(right_65_write_write_en),
      .clk(clk),
      .out(right_65_write_out),
      .done(right_65_write_done)
  );
  
  std_reg #(32) left_65_read (
      .in(left_65_read_in),
      .write_en(left_65_read_write_en),
      .clk(clk),
      .out(left_65_read_out),
      .done(left_65_read_done)
  );
  
  std_reg #(32) top_65_read (
      .in(top_65_read_in),
      .write_en(top_65_read_write_en),
      .clk(clk),
      .out(top_65_read_out),
      .done(top_65_read_done)
  );
  
  mac_pe #() pe_65 (
      .top(pe_65_top),
      .left(pe_65_left),
      .go(pe_65_go),
      .clk(clk),
      .down(pe_65_down),
      .right(pe_65_right),
      .out(pe_65_out),
      .done(pe_65_done)
  );
  
  std_reg #(32) down_64_write (
      .in(down_64_write_in),
      .write_en(down_64_write_write_en),
      .clk(clk),
      .out(down_64_write_out),
      .done(down_64_write_done)
  );
  
  std_reg #(32) right_64_write (
      .in(right_64_write_in),
      .write_en(right_64_write_write_en),
      .clk(clk),
      .out(right_64_write_out),
      .done(right_64_write_done)
  );
  
  std_reg #(32) left_64_read (
      .in(left_64_read_in),
      .write_en(left_64_read_write_en),
      .clk(clk),
      .out(left_64_read_out),
      .done(left_64_read_done)
  );
  
  std_reg #(32) top_64_read (
      .in(top_64_read_in),
      .write_en(top_64_read_write_en),
      .clk(clk),
      .out(top_64_read_out),
      .done(top_64_read_done)
  );
  
  mac_pe #() pe_64 (
      .top(pe_64_top),
      .left(pe_64_left),
      .go(pe_64_go),
      .clk(clk),
      .down(pe_64_down),
      .right(pe_64_right),
      .out(pe_64_out),
      .done(pe_64_done)
  );
  
  std_reg #(32) down_63_write (
      .in(down_63_write_in),
      .write_en(down_63_write_write_en),
      .clk(clk),
      .out(down_63_write_out),
      .done(down_63_write_done)
  );
  
  std_reg #(32) right_63_write (
      .in(right_63_write_in),
      .write_en(right_63_write_write_en),
      .clk(clk),
      .out(right_63_write_out),
      .done(right_63_write_done)
  );
  
  std_reg #(32) left_63_read (
      .in(left_63_read_in),
      .write_en(left_63_read_write_en),
      .clk(clk),
      .out(left_63_read_out),
      .done(left_63_read_done)
  );
  
  std_reg #(32) top_63_read (
      .in(top_63_read_in),
      .write_en(top_63_read_write_en),
      .clk(clk),
      .out(top_63_read_out),
      .done(top_63_read_done)
  );
  
  mac_pe #() pe_63 (
      .top(pe_63_top),
      .left(pe_63_left),
      .go(pe_63_go),
      .clk(clk),
      .down(pe_63_down),
      .right(pe_63_right),
      .out(pe_63_out),
      .done(pe_63_done)
  );
  
  std_reg #(32) down_62_write (
      .in(down_62_write_in),
      .write_en(down_62_write_write_en),
      .clk(clk),
      .out(down_62_write_out),
      .done(down_62_write_done)
  );
  
  std_reg #(32) right_62_write (
      .in(right_62_write_in),
      .write_en(right_62_write_write_en),
      .clk(clk),
      .out(right_62_write_out),
      .done(right_62_write_done)
  );
  
  std_reg #(32) left_62_read (
      .in(left_62_read_in),
      .write_en(left_62_read_write_en),
      .clk(clk),
      .out(left_62_read_out),
      .done(left_62_read_done)
  );
  
  std_reg #(32) top_62_read (
      .in(top_62_read_in),
      .write_en(top_62_read_write_en),
      .clk(clk),
      .out(top_62_read_out),
      .done(top_62_read_done)
  );
  
  mac_pe #() pe_62 (
      .top(pe_62_top),
      .left(pe_62_left),
      .go(pe_62_go),
      .clk(clk),
      .down(pe_62_down),
      .right(pe_62_right),
      .out(pe_62_out),
      .done(pe_62_done)
  );
  
  std_reg #(32) down_61_write (
      .in(down_61_write_in),
      .write_en(down_61_write_write_en),
      .clk(clk),
      .out(down_61_write_out),
      .done(down_61_write_done)
  );
  
  std_reg #(32) right_61_write (
      .in(right_61_write_in),
      .write_en(right_61_write_write_en),
      .clk(clk),
      .out(right_61_write_out),
      .done(right_61_write_done)
  );
  
  std_reg #(32) left_61_read (
      .in(left_61_read_in),
      .write_en(left_61_read_write_en),
      .clk(clk),
      .out(left_61_read_out),
      .done(left_61_read_done)
  );
  
  std_reg #(32) top_61_read (
      .in(top_61_read_in),
      .write_en(top_61_read_write_en),
      .clk(clk),
      .out(top_61_read_out),
      .done(top_61_read_done)
  );
  
  mac_pe #() pe_61 (
      .top(pe_61_top),
      .left(pe_61_left),
      .go(pe_61_go),
      .clk(clk),
      .down(pe_61_down),
      .right(pe_61_right),
      .out(pe_61_out),
      .done(pe_61_done)
  );
  
  std_reg #(32) down_60_write (
      .in(down_60_write_in),
      .write_en(down_60_write_write_en),
      .clk(clk),
      .out(down_60_write_out),
      .done(down_60_write_done)
  );
  
  std_reg #(32) right_60_write (
      .in(right_60_write_in),
      .write_en(right_60_write_write_en),
      .clk(clk),
      .out(right_60_write_out),
      .done(right_60_write_done)
  );
  
  std_reg #(32) left_60_read (
      .in(left_60_read_in),
      .write_en(left_60_read_write_en),
      .clk(clk),
      .out(left_60_read_out),
      .done(left_60_read_done)
  );
  
  std_reg #(32) top_60_read (
      .in(top_60_read_in),
      .write_en(top_60_read_write_en),
      .clk(clk),
      .out(top_60_read_out),
      .done(top_60_read_done)
  );
  
  mac_pe #() pe_60 (
      .top(pe_60_top),
      .left(pe_60_left),
      .go(pe_60_go),
      .clk(clk),
      .down(pe_60_down),
      .right(pe_60_right),
      .out(pe_60_out),
      .done(pe_60_done)
  );
  
  std_reg #(32) down_57_write (
      .in(down_57_write_in),
      .write_en(down_57_write_write_en),
      .clk(clk),
      .out(down_57_write_out),
      .done(down_57_write_done)
  );
  
  std_reg #(32) left_57_read (
      .in(left_57_read_in),
      .write_en(left_57_read_write_en),
      .clk(clk),
      .out(left_57_read_out),
      .done(left_57_read_done)
  );
  
  std_reg #(32) top_57_read (
      .in(top_57_read_in),
      .write_en(top_57_read_write_en),
      .clk(clk),
      .out(top_57_read_out),
      .done(top_57_read_done)
  );
  
  mac_pe #() pe_57 (
      .top(pe_57_top),
      .left(pe_57_left),
      .go(pe_57_go),
      .clk(clk),
      .down(pe_57_down),
      .right(pe_57_right),
      .out(pe_57_out),
      .done(pe_57_done)
  );
  
  std_reg #(32) down_56_write (
      .in(down_56_write_in),
      .write_en(down_56_write_write_en),
      .clk(clk),
      .out(down_56_write_out),
      .done(down_56_write_done)
  );
  
  std_reg #(32) right_56_write (
      .in(right_56_write_in),
      .write_en(right_56_write_write_en),
      .clk(clk),
      .out(right_56_write_out),
      .done(right_56_write_done)
  );
  
  std_reg #(32) left_56_read (
      .in(left_56_read_in),
      .write_en(left_56_read_write_en),
      .clk(clk),
      .out(left_56_read_out),
      .done(left_56_read_done)
  );
  
  std_reg #(32) top_56_read (
      .in(top_56_read_in),
      .write_en(top_56_read_write_en),
      .clk(clk),
      .out(top_56_read_out),
      .done(top_56_read_done)
  );
  
  mac_pe #() pe_56 (
      .top(pe_56_top),
      .left(pe_56_left),
      .go(pe_56_go),
      .clk(clk),
      .down(pe_56_down),
      .right(pe_56_right),
      .out(pe_56_out),
      .done(pe_56_done)
  );
  
  std_reg #(32) down_55_write (
      .in(down_55_write_in),
      .write_en(down_55_write_write_en),
      .clk(clk),
      .out(down_55_write_out),
      .done(down_55_write_done)
  );
  
  std_reg #(32) right_55_write (
      .in(right_55_write_in),
      .write_en(right_55_write_write_en),
      .clk(clk),
      .out(right_55_write_out),
      .done(right_55_write_done)
  );
  
  std_reg #(32) left_55_read (
      .in(left_55_read_in),
      .write_en(left_55_read_write_en),
      .clk(clk),
      .out(left_55_read_out),
      .done(left_55_read_done)
  );
  
  std_reg #(32) top_55_read (
      .in(top_55_read_in),
      .write_en(top_55_read_write_en),
      .clk(clk),
      .out(top_55_read_out),
      .done(top_55_read_done)
  );
  
  mac_pe #() pe_55 (
      .top(pe_55_top),
      .left(pe_55_left),
      .go(pe_55_go),
      .clk(clk),
      .down(pe_55_down),
      .right(pe_55_right),
      .out(pe_55_out),
      .done(pe_55_done)
  );
  
  std_reg #(32) down_54_write (
      .in(down_54_write_in),
      .write_en(down_54_write_write_en),
      .clk(clk),
      .out(down_54_write_out),
      .done(down_54_write_done)
  );
  
  std_reg #(32) right_54_write (
      .in(right_54_write_in),
      .write_en(right_54_write_write_en),
      .clk(clk),
      .out(right_54_write_out),
      .done(right_54_write_done)
  );
  
  std_reg #(32) left_54_read (
      .in(left_54_read_in),
      .write_en(left_54_read_write_en),
      .clk(clk),
      .out(left_54_read_out),
      .done(left_54_read_done)
  );
  
  std_reg #(32) top_54_read (
      .in(top_54_read_in),
      .write_en(top_54_read_write_en),
      .clk(clk),
      .out(top_54_read_out),
      .done(top_54_read_done)
  );
  
  mac_pe #() pe_54 (
      .top(pe_54_top),
      .left(pe_54_left),
      .go(pe_54_go),
      .clk(clk),
      .down(pe_54_down),
      .right(pe_54_right),
      .out(pe_54_out),
      .done(pe_54_done)
  );
  
  std_reg #(32) down_53_write (
      .in(down_53_write_in),
      .write_en(down_53_write_write_en),
      .clk(clk),
      .out(down_53_write_out),
      .done(down_53_write_done)
  );
  
  std_reg #(32) right_53_write (
      .in(right_53_write_in),
      .write_en(right_53_write_write_en),
      .clk(clk),
      .out(right_53_write_out),
      .done(right_53_write_done)
  );
  
  std_reg #(32) left_53_read (
      .in(left_53_read_in),
      .write_en(left_53_read_write_en),
      .clk(clk),
      .out(left_53_read_out),
      .done(left_53_read_done)
  );
  
  std_reg #(32) top_53_read (
      .in(top_53_read_in),
      .write_en(top_53_read_write_en),
      .clk(clk),
      .out(top_53_read_out),
      .done(top_53_read_done)
  );
  
  mac_pe #() pe_53 (
      .top(pe_53_top),
      .left(pe_53_left),
      .go(pe_53_go),
      .clk(clk),
      .down(pe_53_down),
      .right(pe_53_right),
      .out(pe_53_out),
      .done(pe_53_done)
  );
  
  std_reg #(32) down_52_write (
      .in(down_52_write_in),
      .write_en(down_52_write_write_en),
      .clk(clk),
      .out(down_52_write_out),
      .done(down_52_write_done)
  );
  
  std_reg #(32) right_52_write (
      .in(right_52_write_in),
      .write_en(right_52_write_write_en),
      .clk(clk),
      .out(right_52_write_out),
      .done(right_52_write_done)
  );
  
  std_reg #(32) left_52_read (
      .in(left_52_read_in),
      .write_en(left_52_read_write_en),
      .clk(clk),
      .out(left_52_read_out),
      .done(left_52_read_done)
  );
  
  std_reg #(32) top_52_read (
      .in(top_52_read_in),
      .write_en(top_52_read_write_en),
      .clk(clk),
      .out(top_52_read_out),
      .done(top_52_read_done)
  );
  
  mac_pe #() pe_52 (
      .top(pe_52_top),
      .left(pe_52_left),
      .go(pe_52_go),
      .clk(clk),
      .down(pe_52_down),
      .right(pe_52_right),
      .out(pe_52_out),
      .done(pe_52_done)
  );
  
  std_reg #(32) down_51_write (
      .in(down_51_write_in),
      .write_en(down_51_write_write_en),
      .clk(clk),
      .out(down_51_write_out),
      .done(down_51_write_done)
  );
  
  std_reg #(32) right_51_write (
      .in(right_51_write_in),
      .write_en(right_51_write_write_en),
      .clk(clk),
      .out(right_51_write_out),
      .done(right_51_write_done)
  );
  
  std_reg #(32) left_51_read (
      .in(left_51_read_in),
      .write_en(left_51_read_write_en),
      .clk(clk),
      .out(left_51_read_out),
      .done(left_51_read_done)
  );
  
  std_reg #(32) top_51_read (
      .in(top_51_read_in),
      .write_en(top_51_read_write_en),
      .clk(clk),
      .out(top_51_read_out),
      .done(top_51_read_done)
  );
  
  mac_pe #() pe_51 (
      .top(pe_51_top),
      .left(pe_51_left),
      .go(pe_51_go),
      .clk(clk),
      .down(pe_51_down),
      .right(pe_51_right),
      .out(pe_51_out),
      .done(pe_51_done)
  );
  
  std_reg #(32) down_50_write (
      .in(down_50_write_in),
      .write_en(down_50_write_write_en),
      .clk(clk),
      .out(down_50_write_out),
      .done(down_50_write_done)
  );
  
  std_reg #(32) right_50_write (
      .in(right_50_write_in),
      .write_en(right_50_write_write_en),
      .clk(clk),
      .out(right_50_write_out),
      .done(right_50_write_done)
  );
  
  std_reg #(32) left_50_read (
      .in(left_50_read_in),
      .write_en(left_50_read_write_en),
      .clk(clk),
      .out(left_50_read_out),
      .done(left_50_read_done)
  );
  
  std_reg #(32) top_50_read (
      .in(top_50_read_in),
      .write_en(top_50_read_write_en),
      .clk(clk),
      .out(top_50_read_out),
      .done(top_50_read_done)
  );
  
  mac_pe #() pe_50 (
      .top(pe_50_top),
      .left(pe_50_left),
      .go(pe_50_go),
      .clk(clk),
      .down(pe_50_down),
      .right(pe_50_right),
      .out(pe_50_out),
      .done(pe_50_done)
  );
  
  std_reg #(32) down_47_write (
      .in(down_47_write_in),
      .write_en(down_47_write_write_en),
      .clk(clk),
      .out(down_47_write_out),
      .done(down_47_write_done)
  );
  
  std_reg #(32) left_47_read (
      .in(left_47_read_in),
      .write_en(left_47_read_write_en),
      .clk(clk),
      .out(left_47_read_out),
      .done(left_47_read_done)
  );
  
  std_reg #(32) top_47_read (
      .in(top_47_read_in),
      .write_en(top_47_read_write_en),
      .clk(clk),
      .out(top_47_read_out),
      .done(top_47_read_done)
  );
  
  mac_pe #() pe_47 (
      .top(pe_47_top),
      .left(pe_47_left),
      .go(pe_47_go),
      .clk(clk),
      .down(pe_47_down),
      .right(pe_47_right),
      .out(pe_47_out),
      .done(pe_47_done)
  );
  
  std_reg #(32) down_46_write (
      .in(down_46_write_in),
      .write_en(down_46_write_write_en),
      .clk(clk),
      .out(down_46_write_out),
      .done(down_46_write_done)
  );
  
  std_reg #(32) right_46_write (
      .in(right_46_write_in),
      .write_en(right_46_write_write_en),
      .clk(clk),
      .out(right_46_write_out),
      .done(right_46_write_done)
  );
  
  std_reg #(32) left_46_read (
      .in(left_46_read_in),
      .write_en(left_46_read_write_en),
      .clk(clk),
      .out(left_46_read_out),
      .done(left_46_read_done)
  );
  
  std_reg #(32) top_46_read (
      .in(top_46_read_in),
      .write_en(top_46_read_write_en),
      .clk(clk),
      .out(top_46_read_out),
      .done(top_46_read_done)
  );
  
  mac_pe #() pe_46 (
      .top(pe_46_top),
      .left(pe_46_left),
      .go(pe_46_go),
      .clk(clk),
      .down(pe_46_down),
      .right(pe_46_right),
      .out(pe_46_out),
      .done(pe_46_done)
  );
  
  std_reg #(32) down_45_write (
      .in(down_45_write_in),
      .write_en(down_45_write_write_en),
      .clk(clk),
      .out(down_45_write_out),
      .done(down_45_write_done)
  );
  
  std_reg #(32) right_45_write (
      .in(right_45_write_in),
      .write_en(right_45_write_write_en),
      .clk(clk),
      .out(right_45_write_out),
      .done(right_45_write_done)
  );
  
  std_reg #(32) left_45_read (
      .in(left_45_read_in),
      .write_en(left_45_read_write_en),
      .clk(clk),
      .out(left_45_read_out),
      .done(left_45_read_done)
  );
  
  std_reg #(32) top_45_read (
      .in(top_45_read_in),
      .write_en(top_45_read_write_en),
      .clk(clk),
      .out(top_45_read_out),
      .done(top_45_read_done)
  );
  
  mac_pe #() pe_45 (
      .top(pe_45_top),
      .left(pe_45_left),
      .go(pe_45_go),
      .clk(clk),
      .down(pe_45_down),
      .right(pe_45_right),
      .out(pe_45_out),
      .done(pe_45_done)
  );
  
  std_reg #(32) down_44_write (
      .in(down_44_write_in),
      .write_en(down_44_write_write_en),
      .clk(clk),
      .out(down_44_write_out),
      .done(down_44_write_done)
  );
  
  std_reg #(32) right_44_write (
      .in(right_44_write_in),
      .write_en(right_44_write_write_en),
      .clk(clk),
      .out(right_44_write_out),
      .done(right_44_write_done)
  );
  
  std_reg #(32) left_44_read (
      .in(left_44_read_in),
      .write_en(left_44_read_write_en),
      .clk(clk),
      .out(left_44_read_out),
      .done(left_44_read_done)
  );
  
  std_reg #(32) top_44_read (
      .in(top_44_read_in),
      .write_en(top_44_read_write_en),
      .clk(clk),
      .out(top_44_read_out),
      .done(top_44_read_done)
  );
  
  mac_pe #() pe_44 (
      .top(pe_44_top),
      .left(pe_44_left),
      .go(pe_44_go),
      .clk(clk),
      .down(pe_44_down),
      .right(pe_44_right),
      .out(pe_44_out),
      .done(pe_44_done)
  );
  
  std_reg #(32) down_43_write (
      .in(down_43_write_in),
      .write_en(down_43_write_write_en),
      .clk(clk),
      .out(down_43_write_out),
      .done(down_43_write_done)
  );
  
  std_reg #(32) right_43_write (
      .in(right_43_write_in),
      .write_en(right_43_write_write_en),
      .clk(clk),
      .out(right_43_write_out),
      .done(right_43_write_done)
  );
  
  std_reg #(32) left_43_read (
      .in(left_43_read_in),
      .write_en(left_43_read_write_en),
      .clk(clk),
      .out(left_43_read_out),
      .done(left_43_read_done)
  );
  
  std_reg #(32) top_43_read (
      .in(top_43_read_in),
      .write_en(top_43_read_write_en),
      .clk(clk),
      .out(top_43_read_out),
      .done(top_43_read_done)
  );
  
  mac_pe #() pe_43 (
      .top(pe_43_top),
      .left(pe_43_left),
      .go(pe_43_go),
      .clk(clk),
      .down(pe_43_down),
      .right(pe_43_right),
      .out(pe_43_out),
      .done(pe_43_done)
  );
  
  std_reg #(32) down_42_write (
      .in(down_42_write_in),
      .write_en(down_42_write_write_en),
      .clk(clk),
      .out(down_42_write_out),
      .done(down_42_write_done)
  );
  
  std_reg #(32) right_42_write (
      .in(right_42_write_in),
      .write_en(right_42_write_write_en),
      .clk(clk),
      .out(right_42_write_out),
      .done(right_42_write_done)
  );
  
  std_reg #(32) left_42_read (
      .in(left_42_read_in),
      .write_en(left_42_read_write_en),
      .clk(clk),
      .out(left_42_read_out),
      .done(left_42_read_done)
  );
  
  std_reg #(32) top_42_read (
      .in(top_42_read_in),
      .write_en(top_42_read_write_en),
      .clk(clk),
      .out(top_42_read_out),
      .done(top_42_read_done)
  );
  
  mac_pe #() pe_42 (
      .top(pe_42_top),
      .left(pe_42_left),
      .go(pe_42_go),
      .clk(clk),
      .down(pe_42_down),
      .right(pe_42_right),
      .out(pe_42_out),
      .done(pe_42_done)
  );
  
  std_reg #(32) down_41_write (
      .in(down_41_write_in),
      .write_en(down_41_write_write_en),
      .clk(clk),
      .out(down_41_write_out),
      .done(down_41_write_done)
  );
  
  std_reg #(32) right_41_write (
      .in(right_41_write_in),
      .write_en(right_41_write_write_en),
      .clk(clk),
      .out(right_41_write_out),
      .done(right_41_write_done)
  );
  
  std_reg #(32) left_41_read (
      .in(left_41_read_in),
      .write_en(left_41_read_write_en),
      .clk(clk),
      .out(left_41_read_out),
      .done(left_41_read_done)
  );
  
  std_reg #(32) top_41_read (
      .in(top_41_read_in),
      .write_en(top_41_read_write_en),
      .clk(clk),
      .out(top_41_read_out),
      .done(top_41_read_done)
  );
  
  mac_pe #() pe_41 (
      .top(pe_41_top),
      .left(pe_41_left),
      .go(pe_41_go),
      .clk(clk),
      .down(pe_41_down),
      .right(pe_41_right),
      .out(pe_41_out),
      .done(pe_41_done)
  );
  
  std_reg #(32) down_40_write (
      .in(down_40_write_in),
      .write_en(down_40_write_write_en),
      .clk(clk),
      .out(down_40_write_out),
      .done(down_40_write_done)
  );
  
  std_reg #(32) right_40_write (
      .in(right_40_write_in),
      .write_en(right_40_write_write_en),
      .clk(clk),
      .out(right_40_write_out),
      .done(right_40_write_done)
  );
  
  std_reg #(32) left_40_read (
      .in(left_40_read_in),
      .write_en(left_40_read_write_en),
      .clk(clk),
      .out(left_40_read_out),
      .done(left_40_read_done)
  );
  
  std_reg #(32) top_40_read (
      .in(top_40_read_in),
      .write_en(top_40_read_write_en),
      .clk(clk),
      .out(top_40_read_out),
      .done(top_40_read_done)
  );
  
  mac_pe #() pe_40 (
      .top(pe_40_top),
      .left(pe_40_left),
      .go(pe_40_go),
      .clk(clk),
      .down(pe_40_down),
      .right(pe_40_right),
      .out(pe_40_out),
      .done(pe_40_done)
  );
  
  std_reg #(32) down_37_write (
      .in(down_37_write_in),
      .write_en(down_37_write_write_en),
      .clk(clk),
      .out(down_37_write_out),
      .done(down_37_write_done)
  );
  
  std_reg #(32) left_37_read (
      .in(left_37_read_in),
      .write_en(left_37_read_write_en),
      .clk(clk),
      .out(left_37_read_out),
      .done(left_37_read_done)
  );
  
  std_reg #(32) top_37_read (
      .in(top_37_read_in),
      .write_en(top_37_read_write_en),
      .clk(clk),
      .out(top_37_read_out),
      .done(top_37_read_done)
  );
  
  mac_pe #() pe_37 (
      .top(pe_37_top),
      .left(pe_37_left),
      .go(pe_37_go),
      .clk(clk),
      .down(pe_37_down),
      .right(pe_37_right),
      .out(pe_37_out),
      .done(pe_37_done)
  );
  
  std_reg #(32) down_36_write (
      .in(down_36_write_in),
      .write_en(down_36_write_write_en),
      .clk(clk),
      .out(down_36_write_out),
      .done(down_36_write_done)
  );
  
  std_reg #(32) right_36_write (
      .in(right_36_write_in),
      .write_en(right_36_write_write_en),
      .clk(clk),
      .out(right_36_write_out),
      .done(right_36_write_done)
  );
  
  std_reg #(32) left_36_read (
      .in(left_36_read_in),
      .write_en(left_36_read_write_en),
      .clk(clk),
      .out(left_36_read_out),
      .done(left_36_read_done)
  );
  
  std_reg #(32) top_36_read (
      .in(top_36_read_in),
      .write_en(top_36_read_write_en),
      .clk(clk),
      .out(top_36_read_out),
      .done(top_36_read_done)
  );
  
  mac_pe #() pe_36 (
      .top(pe_36_top),
      .left(pe_36_left),
      .go(pe_36_go),
      .clk(clk),
      .down(pe_36_down),
      .right(pe_36_right),
      .out(pe_36_out),
      .done(pe_36_done)
  );
  
  std_reg #(32) down_35_write (
      .in(down_35_write_in),
      .write_en(down_35_write_write_en),
      .clk(clk),
      .out(down_35_write_out),
      .done(down_35_write_done)
  );
  
  std_reg #(32) right_35_write (
      .in(right_35_write_in),
      .write_en(right_35_write_write_en),
      .clk(clk),
      .out(right_35_write_out),
      .done(right_35_write_done)
  );
  
  std_reg #(32) left_35_read (
      .in(left_35_read_in),
      .write_en(left_35_read_write_en),
      .clk(clk),
      .out(left_35_read_out),
      .done(left_35_read_done)
  );
  
  std_reg #(32) top_35_read (
      .in(top_35_read_in),
      .write_en(top_35_read_write_en),
      .clk(clk),
      .out(top_35_read_out),
      .done(top_35_read_done)
  );
  
  mac_pe #() pe_35 (
      .top(pe_35_top),
      .left(pe_35_left),
      .go(pe_35_go),
      .clk(clk),
      .down(pe_35_down),
      .right(pe_35_right),
      .out(pe_35_out),
      .done(pe_35_done)
  );
  
  std_reg #(32) down_34_write (
      .in(down_34_write_in),
      .write_en(down_34_write_write_en),
      .clk(clk),
      .out(down_34_write_out),
      .done(down_34_write_done)
  );
  
  std_reg #(32) right_34_write (
      .in(right_34_write_in),
      .write_en(right_34_write_write_en),
      .clk(clk),
      .out(right_34_write_out),
      .done(right_34_write_done)
  );
  
  std_reg #(32) left_34_read (
      .in(left_34_read_in),
      .write_en(left_34_read_write_en),
      .clk(clk),
      .out(left_34_read_out),
      .done(left_34_read_done)
  );
  
  std_reg #(32) top_34_read (
      .in(top_34_read_in),
      .write_en(top_34_read_write_en),
      .clk(clk),
      .out(top_34_read_out),
      .done(top_34_read_done)
  );
  
  mac_pe #() pe_34 (
      .top(pe_34_top),
      .left(pe_34_left),
      .go(pe_34_go),
      .clk(clk),
      .down(pe_34_down),
      .right(pe_34_right),
      .out(pe_34_out),
      .done(pe_34_done)
  );
  
  std_reg #(32) down_33_write (
      .in(down_33_write_in),
      .write_en(down_33_write_write_en),
      .clk(clk),
      .out(down_33_write_out),
      .done(down_33_write_done)
  );
  
  std_reg #(32) right_33_write (
      .in(right_33_write_in),
      .write_en(right_33_write_write_en),
      .clk(clk),
      .out(right_33_write_out),
      .done(right_33_write_done)
  );
  
  std_reg #(32) left_33_read (
      .in(left_33_read_in),
      .write_en(left_33_read_write_en),
      .clk(clk),
      .out(left_33_read_out),
      .done(left_33_read_done)
  );
  
  std_reg #(32) top_33_read (
      .in(top_33_read_in),
      .write_en(top_33_read_write_en),
      .clk(clk),
      .out(top_33_read_out),
      .done(top_33_read_done)
  );
  
  mac_pe #() pe_33 (
      .top(pe_33_top),
      .left(pe_33_left),
      .go(pe_33_go),
      .clk(clk),
      .down(pe_33_down),
      .right(pe_33_right),
      .out(pe_33_out),
      .done(pe_33_done)
  );
  
  std_reg #(32) down_32_write (
      .in(down_32_write_in),
      .write_en(down_32_write_write_en),
      .clk(clk),
      .out(down_32_write_out),
      .done(down_32_write_done)
  );
  
  std_reg #(32) right_32_write (
      .in(right_32_write_in),
      .write_en(right_32_write_write_en),
      .clk(clk),
      .out(right_32_write_out),
      .done(right_32_write_done)
  );
  
  std_reg #(32) left_32_read (
      .in(left_32_read_in),
      .write_en(left_32_read_write_en),
      .clk(clk),
      .out(left_32_read_out),
      .done(left_32_read_done)
  );
  
  std_reg #(32) top_32_read (
      .in(top_32_read_in),
      .write_en(top_32_read_write_en),
      .clk(clk),
      .out(top_32_read_out),
      .done(top_32_read_done)
  );
  
  mac_pe #() pe_32 (
      .top(pe_32_top),
      .left(pe_32_left),
      .go(pe_32_go),
      .clk(clk),
      .down(pe_32_down),
      .right(pe_32_right),
      .out(pe_32_out),
      .done(pe_32_done)
  );
  
  std_reg #(32) down_31_write (
      .in(down_31_write_in),
      .write_en(down_31_write_write_en),
      .clk(clk),
      .out(down_31_write_out),
      .done(down_31_write_done)
  );
  
  std_reg #(32) right_31_write (
      .in(right_31_write_in),
      .write_en(right_31_write_write_en),
      .clk(clk),
      .out(right_31_write_out),
      .done(right_31_write_done)
  );
  
  std_reg #(32) left_31_read (
      .in(left_31_read_in),
      .write_en(left_31_read_write_en),
      .clk(clk),
      .out(left_31_read_out),
      .done(left_31_read_done)
  );
  
  std_reg #(32) top_31_read (
      .in(top_31_read_in),
      .write_en(top_31_read_write_en),
      .clk(clk),
      .out(top_31_read_out),
      .done(top_31_read_done)
  );
  
  mac_pe #() pe_31 (
      .top(pe_31_top),
      .left(pe_31_left),
      .go(pe_31_go),
      .clk(clk),
      .down(pe_31_down),
      .right(pe_31_right),
      .out(pe_31_out),
      .done(pe_31_done)
  );
  
  std_reg #(32) down_30_write (
      .in(down_30_write_in),
      .write_en(down_30_write_write_en),
      .clk(clk),
      .out(down_30_write_out),
      .done(down_30_write_done)
  );
  
  std_reg #(32) right_30_write (
      .in(right_30_write_in),
      .write_en(right_30_write_write_en),
      .clk(clk),
      .out(right_30_write_out),
      .done(right_30_write_done)
  );
  
  std_reg #(32) left_30_read (
      .in(left_30_read_in),
      .write_en(left_30_read_write_en),
      .clk(clk),
      .out(left_30_read_out),
      .done(left_30_read_done)
  );
  
  std_reg #(32) top_30_read (
      .in(top_30_read_in),
      .write_en(top_30_read_write_en),
      .clk(clk),
      .out(top_30_read_out),
      .done(top_30_read_done)
  );
  
  mac_pe #() pe_30 (
      .top(pe_30_top),
      .left(pe_30_left),
      .go(pe_30_go),
      .clk(clk),
      .down(pe_30_down),
      .right(pe_30_right),
      .out(pe_30_out),
      .done(pe_30_done)
  );
  
  std_reg #(32) down_27_write (
      .in(down_27_write_in),
      .write_en(down_27_write_write_en),
      .clk(clk),
      .out(down_27_write_out),
      .done(down_27_write_done)
  );
  
  std_reg #(32) left_27_read (
      .in(left_27_read_in),
      .write_en(left_27_read_write_en),
      .clk(clk),
      .out(left_27_read_out),
      .done(left_27_read_done)
  );
  
  std_reg #(32) top_27_read (
      .in(top_27_read_in),
      .write_en(top_27_read_write_en),
      .clk(clk),
      .out(top_27_read_out),
      .done(top_27_read_done)
  );
  
  mac_pe #() pe_27 (
      .top(pe_27_top),
      .left(pe_27_left),
      .go(pe_27_go),
      .clk(clk),
      .down(pe_27_down),
      .right(pe_27_right),
      .out(pe_27_out),
      .done(pe_27_done)
  );
  
  std_reg #(32) down_26_write (
      .in(down_26_write_in),
      .write_en(down_26_write_write_en),
      .clk(clk),
      .out(down_26_write_out),
      .done(down_26_write_done)
  );
  
  std_reg #(32) right_26_write (
      .in(right_26_write_in),
      .write_en(right_26_write_write_en),
      .clk(clk),
      .out(right_26_write_out),
      .done(right_26_write_done)
  );
  
  std_reg #(32) left_26_read (
      .in(left_26_read_in),
      .write_en(left_26_read_write_en),
      .clk(clk),
      .out(left_26_read_out),
      .done(left_26_read_done)
  );
  
  std_reg #(32) top_26_read (
      .in(top_26_read_in),
      .write_en(top_26_read_write_en),
      .clk(clk),
      .out(top_26_read_out),
      .done(top_26_read_done)
  );
  
  mac_pe #() pe_26 (
      .top(pe_26_top),
      .left(pe_26_left),
      .go(pe_26_go),
      .clk(clk),
      .down(pe_26_down),
      .right(pe_26_right),
      .out(pe_26_out),
      .done(pe_26_done)
  );
  
  std_reg #(32) down_25_write (
      .in(down_25_write_in),
      .write_en(down_25_write_write_en),
      .clk(clk),
      .out(down_25_write_out),
      .done(down_25_write_done)
  );
  
  std_reg #(32) right_25_write (
      .in(right_25_write_in),
      .write_en(right_25_write_write_en),
      .clk(clk),
      .out(right_25_write_out),
      .done(right_25_write_done)
  );
  
  std_reg #(32) left_25_read (
      .in(left_25_read_in),
      .write_en(left_25_read_write_en),
      .clk(clk),
      .out(left_25_read_out),
      .done(left_25_read_done)
  );
  
  std_reg #(32) top_25_read (
      .in(top_25_read_in),
      .write_en(top_25_read_write_en),
      .clk(clk),
      .out(top_25_read_out),
      .done(top_25_read_done)
  );
  
  mac_pe #() pe_25 (
      .top(pe_25_top),
      .left(pe_25_left),
      .go(pe_25_go),
      .clk(clk),
      .down(pe_25_down),
      .right(pe_25_right),
      .out(pe_25_out),
      .done(pe_25_done)
  );
  
  std_reg #(32) down_24_write (
      .in(down_24_write_in),
      .write_en(down_24_write_write_en),
      .clk(clk),
      .out(down_24_write_out),
      .done(down_24_write_done)
  );
  
  std_reg #(32) right_24_write (
      .in(right_24_write_in),
      .write_en(right_24_write_write_en),
      .clk(clk),
      .out(right_24_write_out),
      .done(right_24_write_done)
  );
  
  std_reg #(32) left_24_read (
      .in(left_24_read_in),
      .write_en(left_24_read_write_en),
      .clk(clk),
      .out(left_24_read_out),
      .done(left_24_read_done)
  );
  
  std_reg #(32) top_24_read (
      .in(top_24_read_in),
      .write_en(top_24_read_write_en),
      .clk(clk),
      .out(top_24_read_out),
      .done(top_24_read_done)
  );
  
  mac_pe #() pe_24 (
      .top(pe_24_top),
      .left(pe_24_left),
      .go(pe_24_go),
      .clk(clk),
      .down(pe_24_down),
      .right(pe_24_right),
      .out(pe_24_out),
      .done(pe_24_done)
  );
  
  std_reg #(32) down_23_write (
      .in(down_23_write_in),
      .write_en(down_23_write_write_en),
      .clk(clk),
      .out(down_23_write_out),
      .done(down_23_write_done)
  );
  
  std_reg #(32) right_23_write (
      .in(right_23_write_in),
      .write_en(right_23_write_write_en),
      .clk(clk),
      .out(right_23_write_out),
      .done(right_23_write_done)
  );
  
  std_reg #(32) left_23_read (
      .in(left_23_read_in),
      .write_en(left_23_read_write_en),
      .clk(clk),
      .out(left_23_read_out),
      .done(left_23_read_done)
  );
  
  std_reg #(32) top_23_read (
      .in(top_23_read_in),
      .write_en(top_23_read_write_en),
      .clk(clk),
      .out(top_23_read_out),
      .done(top_23_read_done)
  );
  
  mac_pe #() pe_23 (
      .top(pe_23_top),
      .left(pe_23_left),
      .go(pe_23_go),
      .clk(clk),
      .down(pe_23_down),
      .right(pe_23_right),
      .out(pe_23_out),
      .done(pe_23_done)
  );
  
  std_reg #(32) down_22_write (
      .in(down_22_write_in),
      .write_en(down_22_write_write_en),
      .clk(clk),
      .out(down_22_write_out),
      .done(down_22_write_done)
  );
  
  std_reg #(32) right_22_write (
      .in(right_22_write_in),
      .write_en(right_22_write_write_en),
      .clk(clk),
      .out(right_22_write_out),
      .done(right_22_write_done)
  );
  
  std_reg #(32) left_22_read (
      .in(left_22_read_in),
      .write_en(left_22_read_write_en),
      .clk(clk),
      .out(left_22_read_out),
      .done(left_22_read_done)
  );
  
  std_reg #(32) top_22_read (
      .in(top_22_read_in),
      .write_en(top_22_read_write_en),
      .clk(clk),
      .out(top_22_read_out),
      .done(top_22_read_done)
  );
  
  mac_pe #() pe_22 (
      .top(pe_22_top),
      .left(pe_22_left),
      .go(pe_22_go),
      .clk(clk),
      .down(pe_22_down),
      .right(pe_22_right),
      .out(pe_22_out),
      .done(pe_22_done)
  );
  
  std_reg #(32) down_21_write (
      .in(down_21_write_in),
      .write_en(down_21_write_write_en),
      .clk(clk),
      .out(down_21_write_out),
      .done(down_21_write_done)
  );
  
  std_reg #(32) right_21_write (
      .in(right_21_write_in),
      .write_en(right_21_write_write_en),
      .clk(clk),
      .out(right_21_write_out),
      .done(right_21_write_done)
  );
  
  std_reg #(32) left_21_read (
      .in(left_21_read_in),
      .write_en(left_21_read_write_en),
      .clk(clk),
      .out(left_21_read_out),
      .done(left_21_read_done)
  );
  
  std_reg #(32) top_21_read (
      .in(top_21_read_in),
      .write_en(top_21_read_write_en),
      .clk(clk),
      .out(top_21_read_out),
      .done(top_21_read_done)
  );
  
  mac_pe #() pe_21 (
      .top(pe_21_top),
      .left(pe_21_left),
      .go(pe_21_go),
      .clk(clk),
      .down(pe_21_down),
      .right(pe_21_right),
      .out(pe_21_out),
      .done(pe_21_done)
  );
  
  std_reg #(32) down_20_write (
      .in(down_20_write_in),
      .write_en(down_20_write_write_en),
      .clk(clk),
      .out(down_20_write_out),
      .done(down_20_write_done)
  );
  
  std_reg #(32) right_20_write (
      .in(right_20_write_in),
      .write_en(right_20_write_write_en),
      .clk(clk),
      .out(right_20_write_out),
      .done(right_20_write_done)
  );
  
  std_reg #(32) left_20_read (
      .in(left_20_read_in),
      .write_en(left_20_read_write_en),
      .clk(clk),
      .out(left_20_read_out),
      .done(left_20_read_done)
  );
  
  std_reg #(32) top_20_read (
      .in(top_20_read_in),
      .write_en(top_20_read_write_en),
      .clk(clk),
      .out(top_20_read_out),
      .done(top_20_read_done)
  );
  
  mac_pe #() pe_20 (
      .top(pe_20_top),
      .left(pe_20_left),
      .go(pe_20_go),
      .clk(clk),
      .down(pe_20_down),
      .right(pe_20_right),
      .out(pe_20_out),
      .done(pe_20_done)
  );
  
  std_reg #(32) down_17_write (
      .in(down_17_write_in),
      .write_en(down_17_write_write_en),
      .clk(clk),
      .out(down_17_write_out),
      .done(down_17_write_done)
  );
  
  std_reg #(32) left_17_read (
      .in(left_17_read_in),
      .write_en(left_17_read_write_en),
      .clk(clk),
      .out(left_17_read_out),
      .done(left_17_read_done)
  );
  
  std_reg #(32) top_17_read (
      .in(top_17_read_in),
      .write_en(top_17_read_write_en),
      .clk(clk),
      .out(top_17_read_out),
      .done(top_17_read_done)
  );
  
  mac_pe #() pe_17 (
      .top(pe_17_top),
      .left(pe_17_left),
      .go(pe_17_go),
      .clk(clk),
      .down(pe_17_down),
      .right(pe_17_right),
      .out(pe_17_out),
      .done(pe_17_done)
  );
  
  std_reg #(32) down_16_write (
      .in(down_16_write_in),
      .write_en(down_16_write_write_en),
      .clk(clk),
      .out(down_16_write_out),
      .done(down_16_write_done)
  );
  
  std_reg #(32) right_16_write (
      .in(right_16_write_in),
      .write_en(right_16_write_write_en),
      .clk(clk),
      .out(right_16_write_out),
      .done(right_16_write_done)
  );
  
  std_reg #(32) left_16_read (
      .in(left_16_read_in),
      .write_en(left_16_read_write_en),
      .clk(clk),
      .out(left_16_read_out),
      .done(left_16_read_done)
  );
  
  std_reg #(32) top_16_read (
      .in(top_16_read_in),
      .write_en(top_16_read_write_en),
      .clk(clk),
      .out(top_16_read_out),
      .done(top_16_read_done)
  );
  
  mac_pe #() pe_16 (
      .top(pe_16_top),
      .left(pe_16_left),
      .go(pe_16_go),
      .clk(clk),
      .down(pe_16_down),
      .right(pe_16_right),
      .out(pe_16_out),
      .done(pe_16_done)
  );
  
  std_reg #(32) down_15_write (
      .in(down_15_write_in),
      .write_en(down_15_write_write_en),
      .clk(clk),
      .out(down_15_write_out),
      .done(down_15_write_done)
  );
  
  std_reg #(32) right_15_write (
      .in(right_15_write_in),
      .write_en(right_15_write_write_en),
      .clk(clk),
      .out(right_15_write_out),
      .done(right_15_write_done)
  );
  
  std_reg #(32) left_15_read (
      .in(left_15_read_in),
      .write_en(left_15_read_write_en),
      .clk(clk),
      .out(left_15_read_out),
      .done(left_15_read_done)
  );
  
  std_reg #(32) top_15_read (
      .in(top_15_read_in),
      .write_en(top_15_read_write_en),
      .clk(clk),
      .out(top_15_read_out),
      .done(top_15_read_done)
  );
  
  mac_pe #() pe_15 (
      .top(pe_15_top),
      .left(pe_15_left),
      .go(pe_15_go),
      .clk(clk),
      .down(pe_15_down),
      .right(pe_15_right),
      .out(pe_15_out),
      .done(pe_15_done)
  );
  
  std_reg #(32) down_14_write (
      .in(down_14_write_in),
      .write_en(down_14_write_write_en),
      .clk(clk),
      .out(down_14_write_out),
      .done(down_14_write_done)
  );
  
  std_reg #(32) right_14_write (
      .in(right_14_write_in),
      .write_en(right_14_write_write_en),
      .clk(clk),
      .out(right_14_write_out),
      .done(right_14_write_done)
  );
  
  std_reg #(32) left_14_read (
      .in(left_14_read_in),
      .write_en(left_14_read_write_en),
      .clk(clk),
      .out(left_14_read_out),
      .done(left_14_read_done)
  );
  
  std_reg #(32) top_14_read (
      .in(top_14_read_in),
      .write_en(top_14_read_write_en),
      .clk(clk),
      .out(top_14_read_out),
      .done(top_14_read_done)
  );
  
  mac_pe #() pe_14 (
      .top(pe_14_top),
      .left(pe_14_left),
      .go(pe_14_go),
      .clk(clk),
      .down(pe_14_down),
      .right(pe_14_right),
      .out(pe_14_out),
      .done(pe_14_done)
  );
  
  std_reg #(32) down_13_write (
      .in(down_13_write_in),
      .write_en(down_13_write_write_en),
      .clk(clk),
      .out(down_13_write_out),
      .done(down_13_write_done)
  );
  
  std_reg #(32) right_13_write (
      .in(right_13_write_in),
      .write_en(right_13_write_write_en),
      .clk(clk),
      .out(right_13_write_out),
      .done(right_13_write_done)
  );
  
  std_reg #(32) left_13_read (
      .in(left_13_read_in),
      .write_en(left_13_read_write_en),
      .clk(clk),
      .out(left_13_read_out),
      .done(left_13_read_done)
  );
  
  std_reg #(32) top_13_read (
      .in(top_13_read_in),
      .write_en(top_13_read_write_en),
      .clk(clk),
      .out(top_13_read_out),
      .done(top_13_read_done)
  );
  
  mac_pe #() pe_13 (
      .top(pe_13_top),
      .left(pe_13_left),
      .go(pe_13_go),
      .clk(clk),
      .down(pe_13_down),
      .right(pe_13_right),
      .out(pe_13_out),
      .done(pe_13_done)
  );
  
  std_reg #(32) down_12_write (
      .in(down_12_write_in),
      .write_en(down_12_write_write_en),
      .clk(clk),
      .out(down_12_write_out),
      .done(down_12_write_done)
  );
  
  std_reg #(32) right_12_write (
      .in(right_12_write_in),
      .write_en(right_12_write_write_en),
      .clk(clk),
      .out(right_12_write_out),
      .done(right_12_write_done)
  );
  
  std_reg #(32) left_12_read (
      .in(left_12_read_in),
      .write_en(left_12_read_write_en),
      .clk(clk),
      .out(left_12_read_out),
      .done(left_12_read_done)
  );
  
  std_reg #(32) top_12_read (
      .in(top_12_read_in),
      .write_en(top_12_read_write_en),
      .clk(clk),
      .out(top_12_read_out),
      .done(top_12_read_done)
  );
  
  mac_pe #() pe_12 (
      .top(pe_12_top),
      .left(pe_12_left),
      .go(pe_12_go),
      .clk(clk),
      .down(pe_12_down),
      .right(pe_12_right),
      .out(pe_12_out),
      .done(pe_12_done)
  );
  
  std_reg #(32) down_11_write (
      .in(down_11_write_in),
      .write_en(down_11_write_write_en),
      .clk(clk),
      .out(down_11_write_out),
      .done(down_11_write_done)
  );
  
  std_reg #(32) right_11_write (
      .in(right_11_write_in),
      .write_en(right_11_write_write_en),
      .clk(clk),
      .out(right_11_write_out),
      .done(right_11_write_done)
  );
  
  std_reg #(32) left_11_read (
      .in(left_11_read_in),
      .write_en(left_11_read_write_en),
      .clk(clk),
      .out(left_11_read_out),
      .done(left_11_read_done)
  );
  
  std_reg #(32) top_11_read (
      .in(top_11_read_in),
      .write_en(top_11_read_write_en),
      .clk(clk),
      .out(top_11_read_out),
      .done(top_11_read_done)
  );
  
  mac_pe #() pe_11 (
      .top(pe_11_top),
      .left(pe_11_left),
      .go(pe_11_go),
      .clk(clk),
      .down(pe_11_down),
      .right(pe_11_right),
      .out(pe_11_out),
      .done(pe_11_done)
  );
  
  std_reg #(32) down_10_write (
      .in(down_10_write_in),
      .write_en(down_10_write_write_en),
      .clk(clk),
      .out(down_10_write_out),
      .done(down_10_write_done)
  );
  
  std_reg #(32) right_10_write (
      .in(right_10_write_in),
      .write_en(right_10_write_write_en),
      .clk(clk),
      .out(right_10_write_out),
      .done(right_10_write_done)
  );
  
  std_reg #(32) left_10_read (
      .in(left_10_read_in),
      .write_en(left_10_read_write_en),
      .clk(clk),
      .out(left_10_read_out),
      .done(left_10_read_done)
  );
  
  std_reg #(32) top_10_read (
      .in(top_10_read_in),
      .write_en(top_10_read_write_en),
      .clk(clk),
      .out(top_10_read_out),
      .done(top_10_read_done)
  );
  
  mac_pe #() pe_10 (
      .top(pe_10_top),
      .left(pe_10_left),
      .go(pe_10_go),
      .clk(clk),
      .down(pe_10_down),
      .right(pe_10_right),
      .out(pe_10_out),
      .done(pe_10_done)
  );
  
  std_reg #(32) down_07_write (
      .in(down_07_write_in),
      .write_en(down_07_write_write_en),
      .clk(clk),
      .out(down_07_write_out),
      .done(down_07_write_done)
  );
  
  std_reg #(32) left_07_read (
      .in(left_07_read_in),
      .write_en(left_07_read_write_en),
      .clk(clk),
      .out(left_07_read_out),
      .done(left_07_read_done)
  );
  
  std_reg #(32) top_07_read (
      .in(top_07_read_in),
      .write_en(top_07_read_write_en),
      .clk(clk),
      .out(top_07_read_out),
      .done(top_07_read_done)
  );
  
  mac_pe #() pe_07 (
      .top(pe_07_top),
      .left(pe_07_left),
      .go(pe_07_go),
      .clk(clk),
      .down(pe_07_down),
      .right(pe_07_right),
      .out(pe_07_out),
      .done(pe_07_done)
  );
  
  std_reg #(32) down_06_write (
      .in(down_06_write_in),
      .write_en(down_06_write_write_en),
      .clk(clk),
      .out(down_06_write_out),
      .done(down_06_write_done)
  );
  
  std_reg #(32) right_06_write (
      .in(right_06_write_in),
      .write_en(right_06_write_write_en),
      .clk(clk),
      .out(right_06_write_out),
      .done(right_06_write_done)
  );
  
  std_reg #(32) left_06_read (
      .in(left_06_read_in),
      .write_en(left_06_read_write_en),
      .clk(clk),
      .out(left_06_read_out),
      .done(left_06_read_done)
  );
  
  std_reg #(32) top_06_read (
      .in(top_06_read_in),
      .write_en(top_06_read_write_en),
      .clk(clk),
      .out(top_06_read_out),
      .done(top_06_read_done)
  );
  
  mac_pe #() pe_06 (
      .top(pe_06_top),
      .left(pe_06_left),
      .go(pe_06_go),
      .clk(clk),
      .down(pe_06_down),
      .right(pe_06_right),
      .out(pe_06_out),
      .done(pe_06_done)
  );
  
  std_reg #(32) down_05_write (
      .in(down_05_write_in),
      .write_en(down_05_write_write_en),
      .clk(clk),
      .out(down_05_write_out),
      .done(down_05_write_done)
  );
  
  std_reg #(32) right_05_write (
      .in(right_05_write_in),
      .write_en(right_05_write_write_en),
      .clk(clk),
      .out(right_05_write_out),
      .done(right_05_write_done)
  );
  
  std_reg #(32) left_05_read (
      .in(left_05_read_in),
      .write_en(left_05_read_write_en),
      .clk(clk),
      .out(left_05_read_out),
      .done(left_05_read_done)
  );
  
  std_reg #(32) top_05_read (
      .in(top_05_read_in),
      .write_en(top_05_read_write_en),
      .clk(clk),
      .out(top_05_read_out),
      .done(top_05_read_done)
  );
  
  mac_pe #() pe_05 (
      .top(pe_05_top),
      .left(pe_05_left),
      .go(pe_05_go),
      .clk(clk),
      .down(pe_05_down),
      .right(pe_05_right),
      .out(pe_05_out),
      .done(pe_05_done)
  );
  
  std_reg #(32) down_04_write (
      .in(down_04_write_in),
      .write_en(down_04_write_write_en),
      .clk(clk),
      .out(down_04_write_out),
      .done(down_04_write_done)
  );
  
  std_reg #(32) right_04_write (
      .in(right_04_write_in),
      .write_en(right_04_write_write_en),
      .clk(clk),
      .out(right_04_write_out),
      .done(right_04_write_done)
  );
  
  std_reg #(32) left_04_read (
      .in(left_04_read_in),
      .write_en(left_04_read_write_en),
      .clk(clk),
      .out(left_04_read_out),
      .done(left_04_read_done)
  );
  
  std_reg #(32) top_04_read (
      .in(top_04_read_in),
      .write_en(top_04_read_write_en),
      .clk(clk),
      .out(top_04_read_out),
      .done(top_04_read_done)
  );
  
  mac_pe #() pe_04 (
      .top(pe_04_top),
      .left(pe_04_left),
      .go(pe_04_go),
      .clk(clk),
      .down(pe_04_down),
      .right(pe_04_right),
      .out(pe_04_out),
      .done(pe_04_done)
  );
  
  std_reg #(32) down_03_write (
      .in(down_03_write_in),
      .write_en(down_03_write_write_en),
      .clk(clk),
      .out(down_03_write_out),
      .done(down_03_write_done)
  );
  
  std_reg #(32) right_03_write (
      .in(right_03_write_in),
      .write_en(right_03_write_write_en),
      .clk(clk),
      .out(right_03_write_out),
      .done(right_03_write_done)
  );
  
  std_reg #(32) left_03_read (
      .in(left_03_read_in),
      .write_en(left_03_read_write_en),
      .clk(clk),
      .out(left_03_read_out),
      .done(left_03_read_done)
  );
  
  std_reg #(32) top_03_read (
      .in(top_03_read_in),
      .write_en(top_03_read_write_en),
      .clk(clk),
      .out(top_03_read_out),
      .done(top_03_read_done)
  );
  
  mac_pe #() pe_03 (
      .top(pe_03_top),
      .left(pe_03_left),
      .go(pe_03_go),
      .clk(clk),
      .down(pe_03_down),
      .right(pe_03_right),
      .out(pe_03_out),
      .done(pe_03_done)
  );
  
  std_reg #(32) down_02_write (
      .in(down_02_write_in),
      .write_en(down_02_write_write_en),
      .clk(clk),
      .out(down_02_write_out),
      .done(down_02_write_done)
  );
  
  std_reg #(32) right_02_write (
      .in(right_02_write_in),
      .write_en(right_02_write_write_en),
      .clk(clk),
      .out(right_02_write_out),
      .done(right_02_write_done)
  );
  
  std_reg #(32) left_02_read (
      .in(left_02_read_in),
      .write_en(left_02_read_write_en),
      .clk(clk),
      .out(left_02_read_out),
      .done(left_02_read_done)
  );
  
  std_reg #(32) top_02_read (
      .in(top_02_read_in),
      .write_en(top_02_read_write_en),
      .clk(clk),
      .out(top_02_read_out),
      .done(top_02_read_done)
  );
  
  mac_pe #() pe_02 (
      .top(pe_02_top),
      .left(pe_02_left),
      .go(pe_02_go),
      .clk(clk),
      .down(pe_02_down),
      .right(pe_02_right),
      .out(pe_02_out),
      .done(pe_02_done)
  );
  
  std_reg #(32) down_01_write (
      .in(down_01_write_in),
      .write_en(down_01_write_write_en),
      .clk(clk),
      .out(down_01_write_out),
      .done(down_01_write_done)
  );
  
  std_reg #(32) right_01_write (
      .in(right_01_write_in),
      .write_en(right_01_write_write_en),
      .clk(clk),
      .out(right_01_write_out),
      .done(right_01_write_done)
  );
  
  std_reg #(32) left_01_read (
      .in(left_01_read_in),
      .write_en(left_01_read_write_en),
      .clk(clk),
      .out(left_01_read_out),
      .done(left_01_read_done)
  );
  
  std_reg #(32) top_01_read (
      .in(top_01_read_in),
      .write_en(top_01_read_write_en),
      .clk(clk),
      .out(top_01_read_out),
      .done(top_01_read_done)
  );
  
  mac_pe #() pe_01 (
      .top(pe_01_top),
      .left(pe_01_left),
      .go(pe_01_go),
      .clk(clk),
      .down(pe_01_down),
      .right(pe_01_right),
      .out(pe_01_out),
      .done(pe_01_done)
  );
  
  std_reg #(32) down_00_write (
      .in(down_00_write_in),
      .write_en(down_00_write_write_en),
      .clk(clk),
      .out(down_00_write_out),
      .done(down_00_write_done)
  );
  
  std_reg #(32) right_00_write (
      .in(right_00_write_in),
      .write_en(right_00_write_write_en),
      .clk(clk),
      .out(right_00_write_out),
      .done(right_00_write_done)
  );
  
  std_reg #(32) left_00_read (
      .in(left_00_read_in),
      .write_en(left_00_read_write_en),
      .clk(clk),
      .out(left_00_read_out),
      .done(left_00_read_done)
  );
  
  std_reg #(32) top_00_read (
      .in(top_00_read_in),
      .write_en(top_00_read_write_en),
      .clk(clk),
      .out(top_00_read_out),
      .done(top_00_read_done)
  );
  
  mac_pe #() pe_00 (
      .top(pe_00_top),
      .left(pe_00_left),
      .go(pe_00_go),
      .clk(clk),
      .down(pe_00_down),
      .right(pe_00_right),
      .out(pe_00_out),
      .done(pe_00_done)
  );
  
  std_mem_d1 #(32, 8, 4) l7 (
      .addr0(l7_addr0),
      .write_data(l7_write_data),
      .write_en(l7_write_en),
      .clk(clk),
      .read_data(l7_read_data),
      .done(l7_done)
  );
  
  std_add #(4) l7_add (
      .left(l7_add_left),
      .right(l7_add_right),
      .out(l7_add_out)
  );
  
  std_reg #(4) l7_idx (
      .in(l7_idx_in),
      .write_en(l7_idx_write_en),
      .clk(clk),
      .out(l7_idx_out),
      .done(l7_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l6 (
      .addr0(l6_addr0),
      .write_data(l6_write_data),
      .write_en(l6_write_en),
      .clk(clk),
      .read_data(l6_read_data),
      .done(l6_done)
  );
  
  std_add #(4) l6_add (
      .left(l6_add_left),
      .right(l6_add_right),
      .out(l6_add_out)
  );
  
  std_reg #(4) l6_idx (
      .in(l6_idx_in),
      .write_en(l6_idx_write_en),
      .clk(clk),
      .out(l6_idx_out),
      .done(l6_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l5 (
      .addr0(l5_addr0),
      .write_data(l5_write_data),
      .write_en(l5_write_en),
      .clk(clk),
      .read_data(l5_read_data),
      .done(l5_done)
  );
  
  std_add #(4) l5_add (
      .left(l5_add_left),
      .right(l5_add_right),
      .out(l5_add_out)
  );
  
  std_reg #(4) l5_idx (
      .in(l5_idx_in),
      .write_en(l5_idx_write_en),
      .clk(clk),
      .out(l5_idx_out),
      .done(l5_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l4 (
      .addr0(l4_addr0),
      .write_data(l4_write_data),
      .write_en(l4_write_en),
      .clk(clk),
      .read_data(l4_read_data),
      .done(l4_done)
  );
  
  std_add #(4) l4_add (
      .left(l4_add_left),
      .right(l4_add_right),
      .out(l4_add_out)
  );
  
  std_reg #(4) l4_idx (
      .in(l4_idx_in),
      .write_en(l4_idx_write_en),
      .clk(clk),
      .out(l4_idx_out),
      .done(l4_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l3 (
      .addr0(l3_addr0),
      .write_data(l3_write_data),
      .write_en(l3_write_en),
      .clk(clk),
      .read_data(l3_read_data),
      .done(l3_done)
  );
  
  std_add #(4) l3_add (
      .left(l3_add_left),
      .right(l3_add_right),
      .out(l3_add_out)
  );
  
  std_reg #(4) l3_idx (
      .in(l3_idx_in),
      .write_en(l3_idx_write_en),
      .clk(clk),
      .out(l3_idx_out),
      .done(l3_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l2 (
      .addr0(l2_addr0),
      .write_data(l2_write_data),
      .write_en(l2_write_en),
      .clk(clk),
      .read_data(l2_read_data),
      .done(l2_done)
  );
  
  std_add #(4) l2_add (
      .left(l2_add_left),
      .right(l2_add_right),
      .out(l2_add_out)
  );
  
  std_reg #(4) l2_idx (
      .in(l2_idx_in),
      .write_en(l2_idx_write_en),
      .clk(clk),
      .out(l2_idx_out),
      .done(l2_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l1 (
      .addr0(l1_addr0),
      .write_data(l1_write_data),
      .write_en(l1_write_en),
      .clk(clk),
      .read_data(l1_read_data),
      .done(l1_done)
  );
  
  std_add #(4) l1_add (
      .left(l1_add_left),
      .right(l1_add_right),
      .out(l1_add_out)
  );
  
  std_reg #(4) l1_idx (
      .in(l1_idx_in),
      .write_en(l1_idx_write_en),
      .clk(clk),
      .out(l1_idx_out),
      .done(l1_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) l0 (
      .addr0(l0_addr0),
      .write_data(l0_write_data),
      .write_en(l0_write_en),
      .clk(clk),
      .read_data(l0_read_data),
      .done(l0_done)
  );
  
  std_add #(4) l0_add (
      .left(l0_add_left),
      .right(l0_add_right),
      .out(l0_add_out)
  );
  
  std_reg #(4) l0_idx (
      .in(l0_idx_in),
      .write_en(l0_idx_write_en),
      .clk(clk),
      .out(l0_idx_out),
      .done(l0_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t7 (
      .addr0(t7_addr0),
      .write_data(t7_write_data),
      .write_en(t7_write_en),
      .clk(clk),
      .read_data(t7_read_data),
      .done(t7_done)
  );
  
  std_add #(4) t7_add (
      .left(t7_add_left),
      .right(t7_add_right),
      .out(t7_add_out)
  );
  
  std_reg #(4) t7_idx (
      .in(t7_idx_in),
      .write_en(t7_idx_write_en),
      .clk(clk),
      .out(t7_idx_out),
      .done(t7_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t6 (
      .addr0(t6_addr0),
      .write_data(t6_write_data),
      .write_en(t6_write_en),
      .clk(clk),
      .read_data(t6_read_data),
      .done(t6_done)
  );
  
  std_add #(4) t6_add (
      .left(t6_add_left),
      .right(t6_add_right),
      .out(t6_add_out)
  );
  
  std_reg #(4) t6_idx (
      .in(t6_idx_in),
      .write_en(t6_idx_write_en),
      .clk(clk),
      .out(t6_idx_out),
      .done(t6_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t5 (
      .addr0(t5_addr0),
      .write_data(t5_write_data),
      .write_en(t5_write_en),
      .clk(clk),
      .read_data(t5_read_data),
      .done(t5_done)
  );
  
  std_add #(4) t5_add (
      .left(t5_add_left),
      .right(t5_add_right),
      .out(t5_add_out)
  );
  
  std_reg #(4) t5_idx (
      .in(t5_idx_in),
      .write_en(t5_idx_write_en),
      .clk(clk),
      .out(t5_idx_out),
      .done(t5_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t4 (
      .addr0(t4_addr0),
      .write_data(t4_write_data),
      .write_en(t4_write_en),
      .clk(clk),
      .read_data(t4_read_data),
      .done(t4_done)
  );
  
  std_add #(4) t4_add (
      .left(t4_add_left),
      .right(t4_add_right),
      .out(t4_add_out)
  );
  
  std_reg #(4) t4_idx (
      .in(t4_idx_in),
      .write_en(t4_idx_write_en),
      .clk(clk),
      .out(t4_idx_out),
      .done(t4_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t3 (
      .addr0(t3_addr0),
      .write_data(t3_write_data),
      .write_en(t3_write_en),
      .clk(clk),
      .read_data(t3_read_data),
      .done(t3_done)
  );
  
  std_add #(4) t3_add (
      .left(t3_add_left),
      .right(t3_add_right),
      .out(t3_add_out)
  );
  
  std_reg #(4) t3_idx (
      .in(t3_idx_in),
      .write_en(t3_idx_write_en),
      .clk(clk),
      .out(t3_idx_out),
      .done(t3_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t2 (
      .addr0(t2_addr0),
      .write_data(t2_write_data),
      .write_en(t2_write_en),
      .clk(clk),
      .read_data(t2_read_data),
      .done(t2_done)
  );
  
  std_add #(4) t2_add (
      .left(t2_add_left),
      .right(t2_add_right),
      .out(t2_add_out)
  );
  
  std_reg #(4) t2_idx (
      .in(t2_idx_in),
      .write_en(t2_idx_write_en),
      .clk(clk),
      .out(t2_idx_out),
      .done(t2_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t1 (
      .addr0(t1_addr0),
      .write_data(t1_write_data),
      .write_en(t1_write_en),
      .clk(clk),
      .read_data(t1_read_data),
      .done(t1_done)
  );
  
  std_add #(4) t1_add (
      .left(t1_add_left),
      .right(t1_add_right),
      .out(t1_add_out)
  );
  
  std_reg #(4) t1_idx (
      .in(t1_idx_in),
      .write_en(t1_idx_write_en),
      .clk(clk),
      .out(t1_idx_out),
      .done(t1_idx_done)
  );
  
  std_mem_d1 #(32, 8, 4) t0 (
      .addr0(t0_addr0),
      .write_data(t0_write_data),
      .write_en(t0_write_en),
      .clk(clk),
      .read_data(t0_read_data),
      .done(t0_done)
  );
  
  std_add #(4) t0_add (
      .left(t0_add_left),
      .right(t0_add_right),
      .out(t0_add_out)
  );
  
  std_reg #(4) t0_idx (
      .in(t0_idx_in),
      .write_en(t0_idx_write_en),
      .clk(clk),
      .out(t0_idx_out),
      .done(t0_idx_done)
  );
  
  std_reg #(1) par_reset0 (
      .in(par_reset0_in),
      .write_en(par_reset0_write_en),
      .clk(clk),
      .out(par_reset0_out),
      .done(par_reset0_done)
  );
  
  std_reg #(1) par_done_reg0 (
      .in(par_done_reg0_in),
      .write_en(par_done_reg0_write_en),
      .clk(clk),
      .out(par_done_reg0_out),
      .done(par_done_reg0_done)
  );
  
  std_reg #(1) par_done_reg1 (
      .in(par_done_reg1_in),
      .write_en(par_done_reg1_write_en),
      .clk(clk),
      .out(par_done_reg1_out),
      .done(par_done_reg1_done)
  );
  
  std_reg #(1) par_done_reg2 (
      .in(par_done_reg2_in),
      .write_en(par_done_reg2_write_en),
      .clk(clk),
      .out(par_done_reg2_out),
      .done(par_done_reg2_done)
  );
  
  std_reg #(1) par_done_reg3 (
      .in(par_done_reg3_in),
      .write_en(par_done_reg3_write_en),
      .clk(clk),
      .out(par_done_reg3_out),
      .done(par_done_reg3_done)
  );
  
  std_reg #(1) par_done_reg4 (
      .in(par_done_reg4_in),
      .write_en(par_done_reg4_write_en),
      .clk(clk),
      .out(par_done_reg4_out),
      .done(par_done_reg4_done)
  );
  
  std_reg #(1) par_done_reg5 (
      .in(par_done_reg5_in),
      .write_en(par_done_reg5_write_en),
      .clk(clk),
      .out(par_done_reg5_out),
      .done(par_done_reg5_done)
  );
  
  std_reg #(1) par_done_reg6 (
      .in(par_done_reg6_in),
      .write_en(par_done_reg6_write_en),
      .clk(clk),
      .out(par_done_reg6_out),
      .done(par_done_reg6_done)
  );
  
  std_reg #(1) par_done_reg7 (
      .in(par_done_reg7_in),
      .write_en(par_done_reg7_write_en),
      .clk(clk),
      .out(par_done_reg7_out),
      .done(par_done_reg7_done)
  );
  
  std_reg #(1) par_done_reg8 (
      .in(par_done_reg8_in),
      .write_en(par_done_reg8_write_en),
      .clk(clk),
      .out(par_done_reg8_out),
      .done(par_done_reg8_done)
  );
  
  std_reg #(1) par_done_reg9 (
      .in(par_done_reg9_in),
      .write_en(par_done_reg9_write_en),
      .clk(clk),
      .out(par_done_reg9_out),
      .done(par_done_reg9_done)
  );
  
  std_reg #(1) par_done_reg10 (
      .in(par_done_reg10_in),
      .write_en(par_done_reg10_write_en),
      .clk(clk),
      .out(par_done_reg10_out),
      .done(par_done_reg10_done)
  );
  
  std_reg #(1) par_done_reg11 (
      .in(par_done_reg11_in),
      .write_en(par_done_reg11_write_en),
      .clk(clk),
      .out(par_done_reg11_out),
      .done(par_done_reg11_done)
  );
  
  std_reg #(1) par_done_reg12 (
      .in(par_done_reg12_in),
      .write_en(par_done_reg12_write_en),
      .clk(clk),
      .out(par_done_reg12_out),
      .done(par_done_reg12_done)
  );
  
  std_reg #(1) par_done_reg13 (
      .in(par_done_reg13_in),
      .write_en(par_done_reg13_write_en),
      .clk(clk),
      .out(par_done_reg13_out),
      .done(par_done_reg13_done)
  );
  
  std_reg #(1) par_done_reg14 (
      .in(par_done_reg14_in),
      .write_en(par_done_reg14_write_en),
      .clk(clk),
      .out(par_done_reg14_out),
      .done(par_done_reg14_done)
  );
  
  std_reg #(1) par_done_reg15 (
      .in(par_done_reg15_in),
      .write_en(par_done_reg15_write_en),
      .clk(clk),
      .out(par_done_reg15_out),
      .done(par_done_reg15_done)
  );
  
  std_reg #(1) par_reset1 (
      .in(par_reset1_in),
      .write_en(par_reset1_write_en),
      .clk(clk),
      .out(par_reset1_out),
      .done(par_reset1_done)
  );
  
  std_reg #(1) par_done_reg16 (
      .in(par_done_reg16_in),
      .write_en(par_done_reg16_write_en),
      .clk(clk),
      .out(par_done_reg16_out),
      .done(par_done_reg16_done)
  );
  
  std_reg #(1) par_done_reg17 (
      .in(par_done_reg17_in),
      .write_en(par_done_reg17_write_en),
      .clk(clk),
      .out(par_done_reg17_out),
      .done(par_done_reg17_done)
  );
  
  std_reg #(1) par_reset2 (
      .in(par_reset2_in),
      .write_en(par_reset2_write_en),
      .clk(clk),
      .out(par_reset2_out),
      .done(par_reset2_done)
  );
  
  std_reg #(1) par_done_reg18 (
      .in(par_done_reg18_in),
      .write_en(par_done_reg18_write_en),
      .clk(clk),
      .out(par_done_reg18_out),
      .done(par_done_reg18_done)
  );
  
  std_reg #(1) par_done_reg19 (
      .in(par_done_reg19_in),
      .write_en(par_done_reg19_write_en),
      .clk(clk),
      .out(par_done_reg19_out),
      .done(par_done_reg19_done)
  );
  
  std_reg #(1) par_reset3 (
      .in(par_reset3_in),
      .write_en(par_reset3_write_en),
      .clk(clk),
      .out(par_reset3_out),
      .done(par_reset3_done)
  );
  
  std_reg #(1) par_done_reg20 (
      .in(par_done_reg20_in),
      .write_en(par_done_reg20_write_en),
      .clk(clk),
      .out(par_done_reg20_out),
      .done(par_done_reg20_done)
  );
  
  std_reg #(1) par_done_reg21 (
      .in(par_done_reg21_in),
      .write_en(par_done_reg21_write_en),
      .clk(clk),
      .out(par_done_reg21_out),
      .done(par_done_reg21_done)
  );
  
  std_reg #(1) par_done_reg22 (
      .in(par_done_reg22_in),
      .write_en(par_done_reg22_write_en),
      .clk(clk),
      .out(par_done_reg22_out),
      .done(par_done_reg22_done)
  );
  
  std_reg #(1) par_done_reg23 (
      .in(par_done_reg23_in),
      .write_en(par_done_reg23_write_en),
      .clk(clk),
      .out(par_done_reg23_out),
      .done(par_done_reg23_done)
  );
  
  std_reg #(1) par_done_reg24 (
      .in(par_done_reg24_in),
      .write_en(par_done_reg24_write_en),
      .clk(clk),
      .out(par_done_reg24_out),
      .done(par_done_reg24_done)
  );
  
  std_reg #(1) par_reset4 (
      .in(par_reset4_in),
      .write_en(par_reset4_write_en),
      .clk(clk),
      .out(par_reset4_out),
      .done(par_reset4_done)
  );
  
  std_reg #(1) par_done_reg25 (
      .in(par_done_reg25_in),
      .write_en(par_done_reg25_write_en),
      .clk(clk),
      .out(par_done_reg25_out),
      .done(par_done_reg25_done)
  );
  
  std_reg #(1) par_done_reg26 (
      .in(par_done_reg26_in),
      .write_en(par_done_reg26_write_en),
      .clk(clk),
      .out(par_done_reg26_out),
      .done(par_done_reg26_done)
  );
  
  std_reg #(1) par_done_reg27 (
      .in(par_done_reg27_in),
      .write_en(par_done_reg27_write_en),
      .clk(clk),
      .out(par_done_reg27_out),
      .done(par_done_reg27_done)
  );
  
  std_reg #(1) par_done_reg28 (
      .in(par_done_reg28_in),
      .write_en(par_done_reg28_write_en),
      .clk(clk),
      .out(par_done_reg28_out),
      .done(par_done_reg28_done)
  );
  
  std_reg #(1) par_done_reg29 (
      .in(par_done_reg29_in),
      .write_en(par_done_reg29_write_en),
      .clk(clk),
      .out(par_done_reg29_out),
      .done(par_done_reg29_done)
  );
  
  std_reg #(1) par_done_reg30 (
      .in(par_done_reg30_in),
      .write_en(par_done_reg30_write_en),
      .clk(clk),
      .out(par_done_reg30_out),
      .done(par_done_reg30_done)
  );
  
  std_reg #(1) par_reset5 (
      .in(par_reset5_in),
      .write_en(par_reset5_write_en),
      .clk(clk),
      .out(par_reset5_out),
      .done(par_reset5_done)
  );
  
  std_reg #(1) par_done_reg31 (
      .in(par_done_reg31_in),
      .write_en(par_done_reg31_write_en),
      .clk(clk),
      .out(par_done_reg31_out),
      .done(par_done_reg31_done)
  );
  
  std_reg #(1) par_done_reg32 (
      .in(par_done_reg32_in),
      .write_en(par_done_reg32_write_en),
      .clk(clk),
      .out(par_done_reg32_out),
      .done(par_done_reg32_done)
  );
  
  std_reg #(1) par_done_reg33 (
      .in(par_done_reg33_in),
      .write_en(par_done_reg33_write_en),
      .clk(clk),
      .out(par_done_reg33_out),
      .done(par_done_reg33_done)
  );
  
  std_reg #(1) par_done_reg34 (
      .in(par_done_reg34_in),
      .write_en(par_done_reg34_write_en),
      .clk(clk),
      .out(par_done_reg34_out),
      .done(par_done_reg34_done)
  );
  
  std_reg #(1) par_done_reg35 (
      .in(par_done_reg35_in),
      .write_en(par_done_reg35_write_en),
      .clk(clk),
      .out(par_done_reg35_out),
      .done(par_done_reg35_done)
  );
  
  std_reg #(1) par_done_reg36 (
      .in(par_done_reg36_in),
      .write_en(par_done_reg36_write_en),
      .clk(clk),
      .out(par_done_reg36_out),
      .done(par_done_reg36_done)
  );
  
  std_reg #(1) par_done_reg37 (
      .in(par_done_reg37_in),
      .write_en(par_done_reg37_write_en),
      .clk(clk),
      .out(par_done_reg37_out),
      .done(par_done_reg37_done)
  );
  
  std_reg #(1) par_done_reg38 (
      .in(par_done_reg38_in),
      .write_en(par_done_reg38_write_en),
      .clk(clk),
      .out(par_done_reg38_out),
      .done(par_done_reg38_done)
  );
  
  std_reg #(1) par_done_reg39 (
      .in(par_done_reg39_in),
      .write_en(par_done_reg39_write_en),
      .clk(clk),
      .out(par_done_reg39_out),
      .done(par_done_reg39_done)
  );
  
  std_reg #(1) par_reset6 (
      .in(par_reset6_in),
      .write_en(par_reset6_write_en),
      .clk(clk),
      .out(par_reset6_out),
      .done(par_reset6_done)
  );
  
  std_reg #(1) par_done_reg40 (
      .in(par_done_reg40_in),
      .write_en(par_done_reg40_write_en),
      .clk(clk),
      .out(par_done_reg40_out),
      .done(par_done_reg40_done)
  );
  
  std_reg #(1) par_done_reg41 (
      .in(par_done_reg41_in),
      .write_en(par_done_reg41_write_en),
      .clk(clk),
      .out(par_done_reg41_out),
      .done(par_done_reg41_done)
  );
  
  std_reg #(1) par_done_reg42 (
      .in(par_done_reg42_in),
      .write_en(par_done_reg42_write_en),
      .clk(clk),
      .out(par_done_reg42_out),
      .done(par_done_reg42_done)
  );
  
  std_reg #(1) par_done_reg43 (
      .in(par_done_reg43_in),
      .write_en(par_done_reg43_write_en),
      .clk(clk),
      .out(par_done_reg43_out),
      .done(par_done_reg43_done)
  );
  
  std_reg #(1) par_done_reg44 (
      .in(par_done_reg44_in),
      .write_en(par_done_reg44_write_en),
      .clk(clk),
      .out(par_done_reg44_out),
      .done(par_done_reg44_done)
  );
  
  std_reg #(1) par_done_reg45 (
      .in(par_done_reg45_in),
      .write_en(par_done_reg45_write_en),
      .clk(clk),
      .out(par_done_reg45_out),
      .done(par_done_reg45_done)
  );
  
  std_reg #(1) par_done_reg46 (
      .in(par_done_reg46_in),
      .write_en(par_done_reg46_write_en),
      .clk(clk),
      .out(par_done_reg46_out),
      .done(par_done_reg46_done)
  );
  
  std_reg #(1) par_done_reg47 (
      .in(par_done_reg47_in),
      .write_en(par_done_reg47_write_en),
      .clk(clk),
      .out(par_done_reg47_out),
      .done(par_done_reg47_done)
  );
  
  std_reg #(1) par_done_reg48 (
      .in(par_done_reg48_in),
      .write_en(par_done_reg48_write_en),
      .clk(clk),
      .out(par_done_reg48_out),
      .done(par_done_reg48_done)
  );
  
  std_reg #(1) par_done_reg49 (
      .in(par_done_reg49_in),
      .write_en(par_done_reg49_write_en),
      .clk(clk),
      .out(par_done_reg49_out),
      .done(par_done_reg49_done)
  );
  
  std_reg #(1) par_done_reg50 (
      .in(par_done_reg50_in),
      .write_en(par_done_reg50_write_en),
      .clk(clk),
      .out(par_done_reg50_out),
      .done(par_done_reg50_done)
  );
  
  std_reg #(1) par_done_reg51 (
      .in(par_done_reg51_in),
      .write_en(par_done_reg51_write_en),
      .clk(clk),
      .out(par_done_reg51_out),
      .done(par_done_reg51_done)
  );
  
  std_reg #(1) par_reset7 (
      .in(par_reset7_in),
      .write_en(par_reset7_write_en),
      .clk(clk),
      .out(par_reset7_out),
      .done(par_reset7_done)
  );
  
  std_reg #(1) par_done_reg52 (
      .in(par_done_reg52_in),
      .write_en(par_done_reg52_write_en),
      .clk(clk),
      .out(par_done_reg52_out),
      .done(par_done_reg52_done)
  );
  
  std_reg #(1) par_done_reg53 (
      .in(par_done_reg53_in),
      .write_en(par_done_reg53_write_en),
      .clk(clk),
      .out(par_done_reg53_out),
      .done(par_done_reg53_done)
  );
  
  std_reg #(1) par_done_reg54 (
      .in(par_done_reg54_in),
      .write_en(par_done_reg54_write_en),
      .clk(clk),
      .out(par_done_reg54_out),
      .done(par_done_reg54_done)
  );
  
  std_reg #(1) par_done_reg55 (
      .in(par_done_reg55_in),
      .write_en(par_done_reg55_write_en),
      .clk(clk),
      .out(par_done_reg55_out),
      .done(par_done_reg55_done)
  );
  
  std_reg #(1) par_done_reg56 (
      .in(par_done_reg56_in),
      .write_en(par_done_reg56_write_en),
      .clk(clk),
      .out(par_done_reg56_out),
      .done(par_done_reg56_done)
  );
  
  std_reg #(1) par_done_reg57 (
      .in(par_done_reg57_in),
      .write_en(par_done_reg57_write_en),
      .clk(clk),
      .out(par_done_reg57_out),
      .done(par_done_reg57_done)
  );
  
  std_reg #(1) par_done_reg58 (
      .in(par_done_reg58_in),
      .write_en(par_done_reg58_write_en),
      .clk(clk),
      .out(par_done_reg58_out),
      .done(par_done_reg58_done)
  );
  
  std_reg #(1) par_done_reg59 (
      .in(par_done_reg59_in),
      .write_en(par_done_reg59_write_en),
      .clk(clk),
      .out(par_done_reg59_out),
      .done(par_done_reg59_done)
  );
  
  std_reg #(1) par_done_reg60 (
      .in(par_done_reg60_in),
      .write_en(par_done_reg60_write_en),
      .clk(clk),
      .out(par_done_reg60_out),
      .done(par_done_reg60_done)
  );
  
  std_reg #(1) par_done_reg61 (
      .in(par_done_reg61_in),
      .write_en(par_done_reg61_write_en),
      .clk(clk),
      .out(par_done_reg61_out),
      .done(par_done_reg61_done)
  );
  
  std_reg #(1) par_done_reg62 (
      .in(par_done_reg62_in),
      .write_en(par_done_reg62_write_en),
      .clk(clk),
      .out(par_done_reg62_out),
      .done(par_done_reg62_done)
  );
  
  std_reg #(1) par_done_reg63 (
      .in(par_done_reg63_in),
      .write_en(par_done_reg63_write_en),
      .clk(clk),
      .out(par_done_reg63_out),
      .done(par_done_reg63_done)
  );
  
  std_reg #(1) par_done_reg64 (
      .in(par_done_reg64_in),
      .write_en(par_done_reg64_write_en),
      .clk(clk),
      .out(par_done_reg64_out),
      .done(par_done_reg64_done)
  );
  
  std_reg #(1) par_done_reg65 (
      .in(par_done_reg65_in),
      .write_en(par_done_reg65_write_en),
      .clk(clk),
      .out(par_done_reg65_out),
      .done(par_done_reg65_done)
  );
  
  std_reg #(1) par_reset8 (
      .in(par_reset8_in),
      .write_en(par_reset8_write_en),
      .clk(clk),
      .out(par_reset8_out),
      .done(par_reset8_done)
  );
  
  std_reg #(1) par_done_reg66 (
      .in(par_done_reg66_in),
      .write_en(par_done_reg66_write_en),
      .clk(clk),
      .out(par_done_reg66_out),
      .done(par_done_reg66_done)
  );
  
  std_reg #(1) par_done_reg67 (
      .in(par_done_reg67_in),
      .write_en(par_done_reg67_write_en),
      .clk(clk),
      .out(par_done_reg67_out),
      .done(par_done_reg67_done)
  );
  
  std_reg #(1) par_done_reg68 (
      .in(par_done_reg68_in),
      .write_en(par_done_reg68_write_en),
      .clk(clk),
      .out(par_done_reg68_out),
      .done(par_done_reg68_done)
  );
  
  std_reg #(1) par_done_reg69 (
      .in(par_done_reg69_in),
      .write_en(par_done_reg69_write_en),
      .clk(clk),
      .out(par_done_reg69_out),
      .done(par_done_reg69_done)
  );
  
  std_reg #(1) par_done_reg70 (
      .in(par_done_reg70_in),
      .write_en(par_done_reg70_write_en),
      .clk(clk),
      .out(par_done_reg70_out),
      .done(par_done_reg70_done)
  );
  
  std_reg #(1) par_done_reg71 (
      .in(par_done_reg71_in),
      .write_en(par_done_reg71_write_en),
      .clk(clk),
      .out(par_done_reg71_out),
      .done(par_done_reg71_done)
  );
  
  std_reg #(1) par_done_reg72 (
      .in(par_done_reg72_in),
      .write_en(par_done_reg72_write_en),
      .clk(clk),
      .out(par_done_reg72_out),
      .done(par_done_reg72_done)
  );
  
  std_reg #(1) par_done_reg73 (
      .in(par_done_reg73_in),
      .write_en(par_done_reg73_write_en),
      .clk(clk),
      .out(par_done_reg73_out),
      .done(par_done_reg73_done)
  );
  
  std_reg #(1) par_done_reg74 (
      .in(par_done_reg74_in),
      .write_en(par_done_reg74_write_en),
      .clk(clk),
      .out(par_done_reg74_out),
      .done(par_done_reg74_done)
  );
  
  std_reg #(1) par_done_reg75 (
      .in(par_done_reg75_in),
      .write_en(par_done_reg75_write_en),
      .clk(clk),
      .out(par_done_reg75_out),
      .done(par_done_reg75_done)
  );
  
  std_reg #(1) par_done_reg76 (
      .in(par_done_reg76_in),
      .write_en(par_done_reg76_write_en),
      .clk(clk),
      .out(par_done_reg76_out),
      .done(par_done_reg76_done)
  );
  
  std_reg #(1) par_done_reg77 (
      .in(par_done_reg77_in),
      .write_en(par_done_reg77_write_en),
      .clk(clk),
      .out(par_done_reg77_out),
      .done(par_done_reg77_done)
  );
  
  std_reg #(1) par_done_reg78 (
      .in(par_done_reg78_in),
      .write_en(par_done_reg78_write_en),
      .clk(clk),
      .out(par_done_reg78_out),
      .done(par_done_reg78_done)
  );
  
  std_reg #(1) par_done_reg79 (
      .in(par_done_reg79_in),
      .write_en(par_done_reg79_write_en),
      .clk(clk),
      .out(par_done_reg79_out),
      .done(par_done_reg79_done)
  );
  
  std_reg #(1) par_done_reg80 (
      .in(par_done_reg80_in),
      .write_en(par_done_reg80_write_en),
      .clk(clk),
      .out(par_done_reg80_out),
      .done(par_done_reg80_done)
  );
  
  std_reg #(1) par_done_reg81 (
      .in(par_done_reg81_in),
      .write_en(par_done_reg81_write_en),
      .clk(clk),
      .out(par_done_reg81_out),
      .done(par_done_reg81_done)
  );
  
  std_reg #(1) par_done_reg82 (
      .in(par_done_reg82_in),
      .write_en(par_done_reg82_write_en),
      .clk(clk),
      .out(par_done_reg82_out),
      .done(par_done_reg82_done)
  );
  
  std_reg #(1) par_done_reg83 (
      .in(par_done_reg83_in),
      .write_en(par_done_reg83_write_en),
      .clk(clk),
      .out(par_done_reg83_out),
      .done(par_done_reg83_done)
  );
  
  std_reg #(1) par_done_reg84 (
      .in(par_done_reg84_in),
      .write_en(par_done_reg84_write_en),
      .clk(clk),
      .out(par_done_reg84_out),
      .done(par_done_reg84_done)
  );
  
  std_reg #(1) par_done_reg85 (
      .in(par_done_reg85_in),
      .write_en(par_done_reg85_write_en),
      .clk(clk),
      .out(par_done_reg85_out),
      .done(par_done_reg85_done)
  );
  
  std_reg #(1) par_reset9 (
      .in(par_reset9_in),
      .write_en(par_reset9_write_en),
      .clk(clk),
      .out(par_reset9_out),
      .done(par_reset9_done)
  );
  
  std_reg #(1) par_done_reg86 (
      .in(par_done_reg86_in),
      .write_en(par_done_reg86_write_en),
      .clk(clk),
      .out(par_done_reg86_out),
      .done(par_done_reg86_done)
  );
  
  std_reg #(1) par_done_reg87 (
      .in(par_done_reg87_in),
      .write_en(par_done_reg87_write_en),
      .clk(clk),
      .out(par_done_reg87_out),
      .done(par_done_reg87_done)
  );
  
  std_reg #(1) par_done_reg88 (
      .in(par_done_reg88_in),
      .write_en(par_done_reg88_write_en),
      .clk(clk),
      .out(par_done_reg88_out),
      .done(par_done_reg88_done)
  );
  
  std_reg #(1) par_done_reg89 (
      .in(par_done_reg89_in),
      .write_en(par_done_reg89_write_en),
      .clk(clk),
      .out(par_done_reg89_out),
      .done(par_done_reg89_done)
  );
  
  std_reg #(1) par_done_reg90 (
      .in(par_done_reg90_in),
      .write_en(par_done_reg90_write_en),
      .clk(clk),
      .out(par_done_reg90_out),
      .done(par_done_reg90_done)
  );
  
  std_reg #(1) par_done_reg91 (
      .in(par_done_reg91_in),
      .write_en(par_done_reg91_write_en),
      .clk(clk),
      .out(par_done_reg91_out),
      .done(par_done_reg91_done)
  );
  
  std_reg #(1) par_done_reg92 (
      .in(par_done_reg92_in),
      .write_en(par_done_reg92_write_en),
      .clk(clk),
      .out(par_done_reg92_out),
      .done(par_done_reg92_done)
  );
  
  std_reg #(1) par_done_reg93 (
      .in(par_done_reg93_in),
      .write_en(par_done_reg93_write_en),
      .clk(clk),
      .out(par_done_reg93_out),
      .done(par_done_reg93_done)
  );
  
  std_reg #(1) par_done_reg94 (
      .in(par_done_reg94_in),
      .write_en(par_done_reg94_write_en),
      .clk(clk),
      .out(par_done_reg94_out),
      .done(par_done_reg94_done)
  );
  
  std_reg #(1) par_done_reg95 (
      .in(par_done_reg95_in),
      .write_en(par_done_reg95_write_en),
      .clk(clk),
      .out(par_done_reg95_out),
      .done(par_done_reg95_done)
  );
  
  std_reg #(1) par_done_reg96 (
      .in(par_done_reg96_in),
      .write_en(par_done_reg96_write_en),
      .clk(clk),
      .out(par_done_reg96_out),
      .done(par_done_reg96_done)
  );
  
  std_reg #(1) par_done_reg97 (
      .in(par_done_reg97_in),
      .write_en(par_done_reg97_write_en),
      .clk(clk),
      .out(par_done_reg97_out),
      .done(par_done_reg97_done)
  );
  
  std_reg #(1) par_done_reg98 (
      .in(par_done_reg98_in),
      .write_en(par_done_reg98_write_en),
      .clk(clk),
      .out(par_done_reg98_out),
      .done(par_done_reg98_done)
  );
  
  std_reg #(1) par_done_reg99 (
      .in(par_done_reg99_in),
      .write_en(par_done_reg99_write_en),
      .clk(clk),
      .out(par_done_reg99_out),
      .done(par_done_reg99_done)
  );
  
  std_reg #(1) par_done_reg100 (
      .in(par_done_reg100_in),
      .write_en(par_done_reg100_write_en),
      .clk(clk),
      .out(par_done_reg100_out),
      .done(par_done_reg100_done)
  );
  
  std_reg #(1) par_done_reg101 (
      .in(par_done_reg101_in),
      .write_en(par_done_reg101_write_en),
      .clk(clk),
      .out(par_done_reg101_out),
      .done(par_done_reg101_done)
  );
  
  std_reg #(1) par_done_reg102 (
      .in(par_done_reg102_in),
      .write_en(par_done_reg102_write_en),
      .clk(clk),
      .out(par_done_reg102_out),
      .done(par_done_reg102_done)
  );
  
  std_reg #(1) par_done_reg103 (
      .in(par_done_reg103_in),
      .write_en(par_done_reg103_write_en),
      .clk(clk),
      .out(par_done_reg103_out),
      .done(par_done_reg103_done)
  );
  
  std_reg #(1) par_done_reg104 (
      .in(par_done_reg104_in),
      .write_en(par_done_reg104_write_en),
      .clk(clk),
      .out(par_done_reg104_out),
      .done(par_done_reg104_done)
  );
  
  std_reg #(1) par_done_reg105 (
      .in(par_done_reg105_in),
      .write_en(par_done_reg105_write_en),
      .clk(clk),
      .out(par_done_reg105_out),
      .done(par_done_reg105_done)
  );
  
  std_reg #(1) par_reset10 (
      .in(par_reset10_in),
      .write_en(par_reset10_write_en),
      .clk(clk),
      .out(par_reset10_out),
      .done(par_reset10_done)
  );
  
  std_reg #(1) par_done_reg106 (
      .in(par_done_reg106_in),
      .write_en(par_done_reg106_write_en),
      .clk(clk),
      .out(par_done_reg106_out),
      .done(par_done_reg106_done)
  );
  
  std_reg #(1) par_done_reg107 (
      .in(par_done_reg107_in),
      .write_en(par_done_reg107_write_en),
      .clk(clk),
      .out(par_done_reg107_out),
      .done(par_done_reg107_done)
  );
  
  std_reg #(1) par_done_reg108 (
      .in(par_done_reg108_in),
      .write_en(par_done_reg108_write_en),
      .clk(clk),
      .out(par_done_reg108_out),
      .done(par_done_reg108_done)
  );
  
  std_reg #(1) par_done_reg109 (
      .in(par_done_reg109_in),
      .write_en(par_done_reg109_write_en),
      .clk(clk),
      .out(par_done_reg109_out),
      .done(par_done_reg109_done)
  );
  
  std_reg #(1) par_done_reg110 (
      .in(par_done_reg110_in),
      .write_en(par_done_reg110_write_en),
      .clk(clk),
      .out(par_done_reg110_out),
      .done(par_done_reg110_done)
  );
  
  std_reg #(1) par_done_reg111 (
      .in(par_done_reg111_in),
      .write_en(par_done_reg111_write_en),
      .clk(clk),
      .out(par_done_reg111_out),
      .done(par_done_reg111_done)
  );
  
  std_reg #(1) par_done_reg112 (
      .in(par_done_reg112_in),
      .write_en(par_done_reg112_write_en),
      .clk(clk),
      .out(par_done_reg112_out),
      .done(par_done_reg112_done)
  );
  
  std_reg #(1) par_done_reg113 (
      .in(par_done_reg113_in),
      .write_en(par_done_reg113_write_en),
      .clk(clk),
      .out(par_done_reg113_out),
      .done(par_done_reg113_done)
  );
  
  std_reg #(1) par_done_reg114 (
      .in(par_done_reg114_in),
      .write_en(par_done_reg114_write_en),
      .clk(clk),
      .out(par_done_reg114_out),
      .done(par_done_reg114_done)
  );
  
  std_reg #(1) par_done_reg115 (
      .in(par_done_reg115_in),
      .write_en(par_done_reg115_write_en),
      .clk(clk),
      .out(par_done_reg115_out),
      .done(par_done_reg115_done)
  );
  
  std_reg #(1) par_done_reg116 (
      .in(par_done_reg116_in),
      .write_en(par_done_reg116_write_en),
      .clk(clk),
      .out(par_done_reg116_out),
      .done(par_done_reg116_done)
  );
  
  std_reg #(1) par_done_reg117 (
      .in(par_done_reg117_in),
      .write_en(par_done_reg117_write_en),
      .clk(clk),
      .out(par_done_reg117_out),
      .done(par_done_reg117_done)
  );
  
  std_reg #(1) par_done_reg118 (
      .in(par_done_reg118_in),
      .write_en(par_done_reg118_write_en),
      .clk(clk),
      .out(par_done_reg118_out),
      .done(par_done_reg118_done)
  );
  
  std_reg #(1) par_done_reg119 (
      .in(par_done_reg119_in),
      .write_en(par_done_reg119_write_en),
      .clk(clk),
      .out(par_done_reg119_out),
      .done(par_done_reg119_done)
  );
  
  std_reg #(1) par_done_reg120 (
      .in(par_done_reg120_in),
      .write_en(par_done_reg120_write_en),
      .clk(clk),
      .out(par_done_reg120_out),
      .done(par_done_reg120_done)
  );
  
  std_reg #(1) par_done_reg121 (
      .in(par_done_reg121_in),
      .write_en(par_done_reg121_write_en),
      .clk(clk),
      .out(par_done_reg121_out),
      .done(par_done_reg121_done)
  );
  
  std_reg #(1) par_done_reg122 (
      .in(par_done_reg122_in),
      .write_en(par_done_reg122_write_en),
      .clk(clk),
      .out(par_done_reg122_out),
      .done(par_done_reg122_done)
  );
  
  std_reg #(1) par_done_reg123 (
      .in(par_done_reg123_in),
      .write_en(par_done_reg123_write_en),
      .clk(clk),
      .out(par_done_reg123_out),
      .done(par_done_reg123_done)
  );
  
  std_reg #(1) par_done_reg124 (
      .in(par_done_reg124_in),
      .write_en(par_done_reg124_write_en),
      .clk(clk),
      .out(par_done_reg124_out),
      .done(par_done_reg124_done)
  );
  
  std_reg #(1) par_done_reg125 (
      .in(par_done_reg125_in),
      .write_en(par_done_reg125_write_en),
      .clk(clk),
      .out(par_done_reg125_out),
      .done(par_done_reg125_done)
  );
  
  std_reg #(1) par_done_reg126 (
      .in(par_done_reg126_in),
      .write_en(par_done_reg126_write_en),
      .clk(clk),
      .out(par_done_reg126_out),
      .done(par_done_reg126_done)
  );
  
  std_reg #(1) par_done_reg127 (
      .in(par_done_reg127_in),
      .write_en(par_done_reg127_write_en),
      .clk(clk),
      .out(par_done_reg127_out),
      .done(par_done_reg127_done)
  );
  
  std_reg #(1) par_done_reg128 (
      .in(par_done_reg128_in),
      .write_en(par_done_reg128_write_en),
      .clk(clk),
      .out(par_done_reg128_out),
      .done(par_done_reg128_done)
  );
  
  std_reg #(1) par_done_reg129 (
      .in(par_done_reg129_in),
      .write_en(par_done_reg129_write_en),
      .clk(clk),
      .out(par_done_reg129_out),
      .done(par_done_reg129_done)
  );
  
  std_reg #(1) par_done_reg130 (
      .in(par_done_reg130_in),
      .write_en(par_done_reg130_write_en),
      .clk(clk),
      .out(par_done_reg130_out),
      .done(par_done_reg130_done)
  );
  
  std_reg #(1) par_done_reg131 (
      .in(par_done_reg131_in),
      .write_en(par_done_reg131_write_en),
      .clk(clk),
      .out(par_done_reg131_out),
      .done(par_done_reg131_done)
  );
  
  std_reg #(1) par_done_reg132 (
      .in(par_done_reg132_in),
      .write_en(par_done_reg132_write_en),
      .clk(clk),
      .out(par_done_reg132_out),
      .done(par_done_reg132_done)
  );
  
  std_reg #(1) par_done_reg133 (
      .in(par_done_reg133_in),
      .write_en(par_done_reg133_write_en),
      .clk(clk),
      .out(par_done_reg133_out),
      .done(par_done_reg133_done)
  );
  
  std_reg #(1) par_done_reg134 (
      .in(par_done_reg134_in),
      .write_en(par_done_reg134_write_en),
      .clk(clk),
      .out(par_done_reg134_out),
      .done(par_done_reg134_done)
  );
  
  std_reg #(1) par_done_reg135 (
      .in(par_done_reg135_in),
      .write_en(par_done_reg135_write_en),
      .clk(clk),
      .out(par_done_reg135_out),
      .done(par_done_reg135_done)
  );
  
  std_reg #(1) par_reset11 (
      .in(par_reset11_in),
      .write_en(par_reset11_write_en),
      .clk(clk),
      .out(par_reset11_out),
      .done(par_reset11_done)
  );
  
  std_reg #(1) par_done_reg136 (
      .in(par_done_reg136_in),
      .write_en(par_done_reg136_write_en),
      .clk(clk),
      .out(par_done_reg136_out),
      .done(par_done_reg136_done)
  );
  
  std_reg #(1) par_done_reg137 (
      .in(par_done_reg137_in),
      .write_en(par_done_reg137_write_en),
      .clk(clk),
      .out(par_done_reg137_out),
      .done(par_done_reg137_done)
  );
  
  std_reg #(1) par_done_reg138 (
      .in(par_done_reg138_in),
      .write_en(par_done_reg138_write_en),
      .clk(clk),
      .out(par_done_reg138_out),
      .done(par_done_reg138_done)
  );
  
  std_reg #(1) par_done_reg139 (
      .in(par_done_reg139_in),
      .write_en(par_done_reg139_write_en),
      .clk(clk),
      .out(par_done_reg139_out),
      .done(par_done_reg139_done)
  );
  
  std_reg #(1) par_done_reg140 (
      .in(par_done_reg140_in),
      .write_en(par_done_reg140_write_en),
      .clk(clk),
      .out(par_done_reg140_out),
      .done(par_done_reg140_done)
  );
  
  std_reg #(1) par_done_reg141 (
      .in(par_done_reg141_in),
      .write_en(par_done_reg141_write_en),
      .clk(clk),
      .out(par_done_reg141_out),
      .done(par_done_reg141_done)
  );
  
  std_reg #(1) par_done_reg142 (
      .in(par_done_reg142_in),
      .write_en(par_done_reg142_write_en),
      .clk(clk),
      .out(par_done_reg142_out),
      .done(par_done_reg142_done)
  );
  
  std_reg #(1) par_done_reg143 (
      .in(par_done_reg143_in),
      .write_en(par_done_reg143_write_en),
      .clk(clk),
      .out(par_done_reg143_out),
      .done(par_done_reg143_done)
  );
  
  std_reg #(1) par_done_reg144 (
      .in(par_done_reg144_in),
      .write_en(par_done_reg144_write_en),
      .clk(clk),
      .out(par_done_reg144_out),
      .done(par_done_reg144_done)
  );
  
  std_reg #(1) par_done_reg145 (
      .in(par_done_reg145_in),
      .write_en(par_done_reg145_write_en),
      .clk(clk),
      .out(par_done_reg145_out),
      .done(par_done_reg145_done)
  );
  
  std_reg #(1) par_done_reg146 (
      .in(par_done_reg146_in),
      .write_en(par_done_reg146_write_en),
      .clk(clk),
      .out(par_done_reg146_out),
      .done(par_done_reg146_done)
  );
  
  std_reg #(1) par_done_reg147 (
      .in(par_done_reg147_in),
      .write_en(par_done_reg147_write_en),
      .clk(clk),
      .out(par_done_reg147_out),
      .done(par_done_reg147_done)
  );
  
  std_reg #(1) par_done_reg148 (
      .in(par_done_reg148_in),
      .write_en(par_done_reg148_write_en),
      .clk(clk),
      .out(par_done_reg148_out),
      .done(par_done_reg148_done)
  );
  
  std_reg #(1) par_done_reg149 (
      .in(par_done_reg149_in),
      .write_en(par_done_reg149_write_en),
      .clk(clk),
      .out(par_done_reg149_out),
      .done(par_done_reg149_done)
  );
  
  std_reg #(1) par_done_reg150 (
      .in(par_done_reg150_in),
      .write_en(par_done_reg150_write_en),
      .clk(clk),
      .out(par_done_reg150_out),
      .done(par_done_reg150_done)
  );
  
  std_reg #(1) par_done_reg151 (
      .in(par_done_reg151_in),
      .write_en(par_done_reg151_write_en),
      .clk(clk),
      .out(par_done_reg151_out),
      .done(par_done_reg151_done)
  );
  
  std_reg #(1) par_done_reg152 (
      .in(par_done_reg152_in),
      .write_en(par_done_reg152_write_en),
      .clk(clk),
      .out(par_done_reg152_out),
      .done(par_done_reg152_done)
  );
  
  std_reg #(1) par_done_reg153 (
      .in(par_done_reg153_in),
      .write_en(par_done_reg153_write_en),
      .clk(clk),
      .out(par_done_reg153_out),
      .done(par_done_reg153_done)
  );
  
  std_reg #(1) par_done_reg154 (
      .in(par_done_reg154_in),
      .write_en(par_done_reg154_write_en),
      .clk(clk),
      .out(par_done_reg154_out),
      .done(par_done_reg154_done)
  );
  
  std_reg #(1) par_done_reg155 (
      .in(par_done_reg155_in),
      .write_en(par_done_reg155_write_en),
      .clk(clk),
      .out(par_done_reg155_out),
      .done(par_done_reg155_done)
  );
  
  std_reg #(1) par_done_reg156 (
      .in(par_done_reg156_in),
      .write_en(par_done_reg156_write_en),
      .clk(clk),
      .out(par_done_reg156_out),
      .done(par_done_reg156_done)
  );
  
  std_reg #(1) par_done_reg157 (
      .in(par_done_reg157_in),
      .write_en(par_done_reg157_write_en),
      .clk(clk),
      .out(par_done_reg157_out),
      .done(par_done_reg157_done)
  );
  
  std_reg #(1) par_done_reg158 (
      .in(par_done_reg158_in),
      .write_en(par_done_reg158_write_en),
      .clk(clk),
      .out(par_done_reg158_out),
      .done(par_done_reg158_done)
  );
  
  std_reg #(1) par_done_reg159 (
      .in(par_done_reg159_in),
      .write_en(par_done_reg159_write_en),
      .clk(clk),
      .out(par_done_reg159_out),
      .done(par_done_reg159_done)
  );
  
  std_reg #(1) par_done_reg160 (
      .in(par_done_reg160_in),
      .write_en(par_done_reg160_write_en),
      .clk(clk),
      .out(par_done_reg160_out),
      .done(par_done_reg160_done)
  );
  
  std_reg #(1) par_done_reg161 (
      .in(par_done_reg161_in),
      .write_en(par_done_reg161_write_en),
      .clk(clk),
      .out(par_done_reg161_out),
      .done(par_done_reg161_done)
  );
  
  std_reg #(1) par_done_reg162 (
      .in(par_done_reg162_in),
      .write_en(par_done_reg162_write_en),
      .clk(clk),
      .out(par_done_reg162_out),
      .done(par_done_reg162_done)
  );
  
  std_reg #(1) par_reset12 (
      .in(par_reset12_in),
      .write_en(par_reset12_write_en),
      .clk(clk),
      .out(par_reset12_out),
      .done(par_reset12_done)
  );
  
  std_reg #(1) par_done_reg163 (
      .in(par_done_reg163_in),
      .write_en(par_done_reg163_write_en),
      .clk(clk),
      .out(par_done_reg163_out),
      .done(par_done_reg163_done)
  );
  
  std_reg #(1) par_done_reg164 (
      .in(par_done_reg164_in),
      .write_en(par_done_reg164_write_en),
      .clk(clk),
      .out(par_done_reg164_out),
      .done(par_done_reg164_done)
  );
  
  std_reg #(1) par_done_reg165 (
      .in(par_done_reg165_in),
      .write_en(par_done_reg165_write_en),
      .clk(clk),
      .out(par_done_reg165_out),
      .done(par_done_reg165_done)
  );
  
  std_reg #(1) par_done_reg166 (
      .in(par_done_reg166_in),
      .write_en(par_done_reg166_write_en),
      .clk(clk),
      .out(par_done_reg166_out),
      .done(par_done_reg166_done)
  );
  
  std_reg #(1) par_done_reg167 (
      .in(par_done_reg167_in),
      .write_en(par_done_reg167_write_en),
      .clk(clk),
      .out(par_done_reg167_out),
      .done(par_done_reg167_done)
  );
  
  std_reg #(1) par_done_reg168 (
      .in(par_done_reg168_in),
      .write_en(par_done_reg168_write_en),
      .clk(clk),
      .out(par_done_reg168_out),
      .done(par_done_reg168_done)
  );
  
  std_reg #(1) par_done_reg169 (
      .in(par_done_reg169_in),
      .write_en(par_done_reg169_write_en),
      .clk(clk),
      .out(par_done_reg169_out),
      .done(par_done_reg169_done)
  );
  
  std_reg #(1) par_done_reg170 (
      .in(par_done_reg170_in),
      .write_en(par_done_reg170_write_en),
      .clk(clk),
      .out(par_done_reg170_out),
      .done(par_done_reg170_done)
  );
  
  std_reg #(1) par_done_reg171 (
      .in(par_done_reg171_in),
      .write_en(par_done_reg171_write_en),
      .clk(clk),
      .out(par_done_reg171_out),
      .done(par_done_reg171_done)
  );
  
  std_reg #(1) par_done_reg172 (
      .in(par_done_reg172_in),
      .write_en(par_done_reg172_write_en),
      .clk(clk),
      .out(par_done_reg172_out),
      .done(par_done_reg172_done)
  );
  
  std_reg #(1) par_done_reg173 (
      .in(par_done_reg173_in),
      .write_en(par_done_reg173_write_en),
      .clk(clk),
      .out(par_done_reg173_out),
      .done(par_done_reg173_done)
  );
  
  std_reg #(1) par_done_reg174 (
      .in(par_done_reg174_in),
      .write_en(par_done_reg174_write_en),
      .clk(clk),
      .out(par_done_reg174_out),
      .done(par_done_reg174_done)
  );
  
  std_reg #(1) par_done_reg175 (
      .in(par_done_reg175_in),
      .write_en(par_done_reg175_write_en),
      .clk(clk),
      .out(par_done_reg175_out),
      .done(par_done_reg175_done)
  );
  
  std_reg #(1) par_done_reg176 (
      .in(par_done_reg176_in),
      .write_en(par_done_reg176_write_en),
      .clk(clk),
      .out(par_done_reg176_out),
      .done(par_done_reg176_done)
  );
  
  std_reg #(1) par_done_reg177 (
      .in(par_done_reg177_in),
      .write_en(par_done_reg177_write_en),
      .clk(clk),
      .out(par_done_reg177_out),
      .done(par_done_reg177_done)
  );
  
  std_reg #(1) par_done_reg178 (
      .in(par_done_reg178_in),
      .write_en(par_done_reg178_write_en),
      .clk(clk),
      .out(par_done_reg178_out),
      .done(par_done_reg178_done)
  );
  
  std_reg #(1) par_done_reg179 (
      .in(par_done_reg179_in),
      .write_en(par_done_reg179_write_en),
      .clk(clk),
      .out(par_done_reg179_out),
      .done(par_done_reg179_done)
  );
  
  std_reg #(1) par_done_reg180 (
      .in(par_done_reg180_in),
      .write_en(par_done_reg180_write_en),
      .clk(clk),
      .out(par_done_reg180_out),
      .done(par_done_reg180_done)
  );
  
  std_reg #(1) par_done_reg181 (
      .in(par_done_reg181_in),
      .write_en(par_done_reg181_write_en),
      .clk(clk),
      .out(par_done_reg181_out),
      .done(par_done_reg181_done)
  );
  
  std_reg #(1) par_done_reg182 (
      .in(par_done_reg182_in),
      .write_en(par_done_reg182_write_en),
      .clk(clk),
      .out(par_done_reg182_out),
      .done(par_done_reg182_done)
  );
  
  std_reg #(1) par_done_reg183 (
      .in(par_done_reg183_in),
      .write_en(par_done_reg183_write_en),
      .clk(clk),
      .out(par_done_reg183_out),
      .done(par_done_reg183_done)
  );
  
  std_reg #(1) par_done_reg184 (
      .in(par_done_reg184_in),
      .write_en(par_done_reg184_write_en),
      .clk(clk),
      .out(par_done_reg184_out),
      .done(par_done_reg184_done)
  );
  
  std_reg #(1) par_done_reg185 (
      .in(par_done_reg185_in),
      .write_en(par_done_reg185_write_en),
      .clk(clk),
      .out(par_done_reg185_out),
      .done(par_done_reg185_done)
  );
  
  std_reg #(1) par_done_reg186 (
      .in(par_done_reg186_in),
      .write_en(par_done_reg186_write_en),
      .clk(clk),
      .out(par_done_reg186_out),
      .done(par_done_reg186_done)
  );
  
  std_reg #(1) par_done_reg187 (
      .in(par_done_reg187_in),
      .write_en(par_done_reg187_write_en),
      .clk(clk),
      .out(par_done_reg187_out),
      .done(par_done_reg187_done)
  );
  
  std_reg #(1) par_done_reg188 (
      .in(par_done_reg188_in),
      .write_en(par_done_reg188_write_en),
      .clk(clk),
      .out(par_done_reg188_out),
      .done(par_done_reg188_done)
  );
  
  std_reg #(1) par_done_reg189 (
      .in(par_done_reg189_in),
      .write_en(par_done_reg189_write_en),
      .clk(clk),
      .out(par_done_reg189_out),
      .done(par_done_reg189_done)
  );
  
  std_reg #(1) par_done_reg190 (
      .in(par_done_reg190_in),
      .write_en(par_done_reg190_write_en),
      .clk(clk),
      .out(par_done_reg190_out),
      .done(par_done_reg190_done)
  );
  
  std_reg #(1) par_done_reg191 (
      .in(par_done_reg191_in),
      .write_en(par_done_reg191_write_en),
      .clk(clk),
      .out(par_done_reg191_out),
      .done(par_done_reg191_done)
  );
  
  std_reg #(1) par_done_reg192 (
      .in(par_done_reg192_in),
      .write_en(par_done_reg192_write_en),
      .clk(clk),
      .out(par_done_reg192_out),
      .done(par_done_reg192_done)
  );
  
  std_reg #(1) par_done_reg193 (
      .in(par_done_reg193_in),
      .write_en(par_done_reg193_write_en),
      .clk(clk),
      .out(par_done_reg193_out),
      .done(par_done_reg193_done)
  );
  
  std_reg #(1) par_done_reg194 (
      .in(par_done_reg194_in),
      .write_en(par_done_reg194_write_en),
      .clk(clk),
      .out(par_done_reg194_out),
      .done(par_done_reg194_done)
  );
  
  std_reg #(1) par_done_reg195 (
      .in(par_done_reg195_in),
      .write_en(par_done_reg195_write_en),
      .clk(clk),
      .out(par_done_reg195_out),
      .done(par_done_reg195_done)
  );
  
  std_reg #(1) par_done_reg196 (
      .in(par_done_reg196_in),
      .write_en(par_done_reg196_write_en),
      .clk(clk),
      .out(par_done_reg196_out),
      .done(par_done_reg196_done)
  );
  
  std_reg #(1) par_done_reg197 (
      .in(par_done_reg197_in),
      .write_en(par_done_reg197_write_en),
      .clk(clk),
      .out(par_done_reg197_out),
      .done(par_done_reg197_done)
  );
  
  std_reg #(1) par_done_reg198 (
      .in(par_done_reg198_in),
      .write_en(par_done_reg198_write_en),
      .clk(clk),
      .out(par_done_reg198_out),
      .done(par_done_reg198_done)
  );
  
  std_reg #(1) par_done_reg199 (
      .in(par_done_reg199_in),
      .write_en(par_done_reg199_write_en),
      .clk(clk),
      .out(par_done_reg199_out),
      .done(par_done_reg199_done)
  );
  
  std_reg #(1) par_done_reg200 (
      .in(par_done_reg200_in),
      .write_en(par_done_reg200_write_en),
      .clk(clk),
      .out(par_done_reg200_out),
      .done(par_done_reg200_done)
  );
  
  std_reg #(1) par_done_reg201 (
      .in(par_done_reg201_in),
      .write_en(par_done_reg201_write_en),
      .clk(clk),
      .out(par_done_reg201_out),
      .done(par_done_reg201_done)
  );
  
  std_reg #(1) par_done_reg202 (
      .in(par_done_reg202_in),
      .write_en(par_done_reg202_write_en),
      .clk(clk),
      .out(par_done_reg202_out),
      .done(par_done_reg202_done)
  );
  
  std_reg #(1) par_done_reg203 (
      .in(par_done_reg203_in),
      .write_en(par_done_reg203_write_en),
      .clk(clk),
      .out(par_done_reg203_out),
      .done(par_done_reg203_done)
  );
  
  std_reg #(1) par_done_reg204 (
      .in(par_done_reg204_in),
      .write_en(par_done_reg204_write_en),
      .clk(clk),
      .out(par_done_reg204_out),
      .done(par_done_reg204_done)
  );
  
  std_reg #(1) par_reset13 (
      .in(par_reset13_in),
      .write_en(par_reset13_write_en),
      .clk(clk),
      .out(par_reset13_out),
      .done(par_reset13_done)
  );
  
  std_reg #(1) par_done_reg205 (
      .in(par_done_reg205_in),
      .write_en(par_done_reg205_write_en),
      .clk(clk),
      .out(par_done_reg205_out),
      .done(par_done_reg205_done)
  );
  
  std_reg #(1) par_done_reg206 (
      .in(par_done_reg206_in),
      .write_en(par_done_reg206_write_en),
      .clk(clk),
      .out(par_done_reg206_out),
      .done(par_done_reg206_done)
  );
  
  std_reg #(1) par_done_reg207 (
      .in(par_done_reg207_in),
      .write_en(par_done_reg207_write_en),
      .clk(clk),
      .out(par_done_reg207_out),
      .done(par_done_reg207_done)
  );
  
  std_reg #(1) par_done_reg208 (
      .in(par_done_reg208_in),
      .write_en(par_done_reg208_write_en),
      .clk(clk),
      .out(par_done_reg208_out),
      .done(par_done_reg208_done)
  );
  
  std_reg #(1) par_done_reg209 (
      .in(par_done_reg209_in),
      .write_en(par_done_reg209_write_en),
      .clk(clk),
      .out(par_done_reg209_out),
      .done(par_done_reg209_done)
  );
  
  std_reg #(1) par_done_reg210 (
      .in(par_done_reg210_in),
      .write_en(par_done_reg210_write_en),
      .clk(clk),
      .out(par_done_reg210_out),
      .done(par_done_reg210_done)
  );
  
  std_reg #(1) par_done_reg211 (
      .in(par_done_reg211_in),
      .write_en(par_done_reg211_write_en),
      .clk(clk),
      .out(par_done_reg211_out),
      .done(par_done_reg211_done)
  );
  
  std_reg #(1) par_done_reg212 (
      .in(par_done_reg212_in),
      .write_en(par_done_reg212_write_en),
      .clk(clk),
      .out(par_done_reg212_out),
      .done(par_done_reg212_done)
  );
  
  std_reg #(1) par_done_reg213 (
      .in(par_done_reg213_in),
      .write_en(par_done_reg213_write_en),
      .clk(clk),
      .out(par_done_reg213_out),
      .done(par_done_reg213_done)
  );
  
  std_reg #(1) par_done_reg214 (
      .in(par_done_reg214_in),
      .write_en(par_done_reg214_write_en),
      .clk(clk),
      .out(par_done_reg214_out),
      .done(par_done_reg214_done)
  );
  
  std_reg #(1) par_done_reg215 (
      .in(par_done_reg215_in),
      .write_en(par_done_reg215_write_en),
      .clk(clk),
      .out(par_done_reg215_out),
      .done(par_done_reg215_done)
  );
  
  std_reg #(1) par_done_reg216 (
      .in(par_done_reg216_in),
      .write_en(par_done_reg216_write_en),
      .clk(clk),
      .out(par_done_reg216_out),
      .done(par_done_reg216_done)
  );
  
  std_reg #(1) par_done_reg217 (
      .in(par_done_reg217_in),
      .write_en(par_done_reg217_write_en),
      .clk(clk),
      .out(par_done_reg217_out),
      .done(par_done_reg217_done)
  );
  
  std_reg #(1) par_done_reg218 (
      .in(par_done_reg218_in),
      .write_en(par_done_reg218_write_en),
      .clk(clk),
      .out(par_done_reg218_out),
      .done(par_done_reg218_done)
  );
  
  std_reg #(1) par_done_reg219 (
      .in(par_done_reg219_in),
      .write_en(par_done_reg219_write_en),
      .clk(clk),
      .out(par_done_reg219_out),
      .done(par_done_reg219_done)
  );
  
  std_reg #(1) par_done_reg220 (
      .in(par_done_reg220_in),
      .write_en(par_done_reg220_write_en),
      .clk(clk),
      .out(par_done_reg220_out),
      .done(par_done_reg220_done)
  );
  
  std_reg #(1) par_done_reg221 (
      .in(par_done_reg221_in),
      .write_en(par_done_reg221_write_en),
      .clk(clk),
      .out(par_done_reg221_out),
      .done(par_done_reg221_done)
  );
  
  std_reg #(1) par_done_reg222 (
      .in(par_done_reg222_in),
      .write_en(par_done_reg222_write_en),
      .clk(clk),
      .out(par_done_reg222_out),
      .done(par_done_reg222_done)
  );
  
  std_reg #(1) par_done_reg223 (
      .in(par_done_reg223_in),
      .write_en(par_done_reg223_write_en),
      .clk(clk),
      .out(par_done_reg223_out),
      .done(par_done_reg223_done)
  );
  
  std_reg #(1) par_done_reg224 (
      .in(par_done_reg224_in),
      .write_en(par_done_reg224_write_en),
      .clk(clk),
      .out(par_done_reg224_out),
      .done(par_done_reg224_done)
  );
  
  std_reg #(1) par_done_reg225 (
      .in(par_done_reg225_in),
      .write_en(par_done_reg225_write_en),
      .clk(clk),
      .out(par_done_reg225_out),
      .done(par_done_reg225_done)
  );
  
  std_reg #(1) par_done_reg226 (
      .in(par_done_reg226_in),
      .write_en(par_done_reg226_write_en),
      .clk(clk),
      .out(par_done_reg226_out),
      .done(par_done_reg226_done)
  );
  
  std_reg #(1) par_done_reg227 (
      .in(par_done_reg227_in),
      .write_en(par_done_reg227_write_en),
      .clk(clk),
      .out(par_done_reg227_out),
      .done(par_done_reg227_done)
  );
  
  std_reg #(1) par_done_reg228 (
      .in(par_done_reg228_in),
      .write_en(par_done_reg228_write_en),
      .clk(clk),
      .out(par_done_reg228_out),
      .done(par_done_reg228_done)
  );
  
  std_reg #(1) par_done_reg229 (
      .in(par_done_reg229_in),
      .write_en(par_done_reg229_write_en),
      .clk(clk),
      .out(par_done_reg229_out),
      .done(par_done_reg229_done)
  );
  
  std_reg #(1) par_done_reg230 (
      .in(par_done_reg230_in),
      .write_en(par_done_reg230_write_en),
      .clk(clk),
      .out(par_done_reg230_out),
      .done(par_done_reg230_done)
  );
  
  std_reg #(1) par_done_reg231 (
      .in(par_done_reg231_in),
      .write_en(par_done_reg231_write_en),
      .clk(clk),
      .out(par_done_reg231_out),
      .done(par_done_reg231_done)
  );
  
  std_reg #(1) par_done_reg232 (
      .in(par_done_reg232_in),
      .write_en(par_done_reg232_write_en),
      .clk(clk),
      .out(par_done_reg232_out),
      .done(par_done_reg232_done)
  );
  
  std_reg #(1) par_done_reg233 (
      .in(par_done_reg233_in),
      .write_en(par_done_reg233_write_en),
      .clk(clk),
      .out(par_done_reg233_out),
      .done(par_done_reg233_done)
  );
  
  std_reg #(1) par_done_reg234 (
      .in(par_done_reg234_in),
      .write_en(par_done_reg234_write_en),
      .clk(clk),
      .out(par_done_reg234_out),
      .done(par_done_reg234_done)
  );
  
  std_reg #(1) par_done_reg235 (
      .in(par_done_reg235_in),
      .write_en(par_done_reg235_write_en),
      .clk(clk),
      .out(par_done_reg235_out),
      .done(par_done_reg235_done)
  );
  
  std_reg #(1) par_done_reg236 (
      .in(par_done_reg236_in),
      .write_en(par_done_reg236_write_en),
      .clk(clk),
      .out(par_done_reg236_out),
      .done(par_done_reg236_done)
  );
  
  std_reg #(1) par_done_reg237 (
      .in(par_done_reg237_in),
      .write_en(par_done_reg237_write_en),
      .clk(clk),
      .out(par_done_reg237_out),
      .done(par_done_reg237_done)
  );
  
  std_reg #(1) par_done_reg238 (
      .in(par_done_reg238_in),
      .write_en(par_done_reg238_write_en),
      .clk(clk),
      .out(par_done_reg238_out),
      .done(par_done_reg238_done)
  );
  
  std_reg #(1) par_done_reg239 (
      .in(par_done_reg239_in),
      .write_en(par_done_reg239_write_en),
      .clk(clk),
      .out(par_done_reg239_out),
      .done(par_done_reg239_done)
  );
  
  std_reg #(1) par_reset14 (
      .in(par_reset14_in),
      .write_en(par_reset14_write_en),
      .clk(clk),
      .out(par_reset14_out),
      .done(par_reset14_done)
  );
  
  std_reg #(1) par_done_reg240 (
      .in(par_done_reg240_in),
      .write_en(par_done_reg240_write_en),
      .clk(clk),
      .out(par_done_reg240_out),
      .done(par_done_reg240_done)
  );
  
  std_reg #(1) par_done_reg241 (
      .in(par_done_reg241_in),
      .write_en(par_done_reg241_write_en),
      .clk(clk),
      .out(par_done_reg241_out),
      .done(par_done_reg241_done)
  );
  
  std_reg #(1) par_done_reg242 (
      .in(par_done_reg242_in),
      .write_en(par_done_reg242_write_en),
      .clk(clk),
      .out(par_done_reg242_out),
      .done(par_done_reg242_done)
  );
  
  std_reg #(1) par_done_reg243 (
      .in(par_done_reg243_in),
      .write_en(par_done_reg243_write_en),
      .clk(clk),
      .out(par_done_reg243_out),
      .done(par_done_reg243_done)
  );
  
  std_reg #(1) par_done_reg244 (
      .in(par_done_reg244_in),
      .write_en(par_done_reg244_write_en),
      .clk(clk),
      .out(par_done_reg244_out),
      .done(par_done_reg244_done)
  );
  
  std_reg #(1) par_done_reg245 (
      .in(par_done_reg245_in),
      .write_en(par_done_reg245_write_en),
      .clk(clk),
      .out(par_done_reg245_out),
      .done(par_done_reg245_done)
  );
  
  std_reg #(1) par_done_reg246 (
      .in(par_done_reg246_in),
      .write_en(par_done_reg246_write_en),
      .clk(clk),
      .out(par_done_reg246_out),
      .done(par_done_reg246_done)
  );
  
  std_reg #(1) par_done_reg247 (
      .in(par_done_reg247_in),
      .write_en(par_done_reg247_write_en),
      .clk(clk),
      .out(par_done_reg247_out),
      .done(par_done_reg247_done)
  );
  
  std_reg #(1) par_done_reg248 (
      .in(par_done_reg248_in),
      .write_en(par_done_reg248_write_en),
      .clk(clk),
      .out(par_done_reg248_out),
      .done(par_done_reg248_done)
  );
  
  std_reg #(1) par_done_reg249 (
      .in(par_done_reg249_in),
      .write_en(par_done_reg249_write_en),
      .clk(clk),
      .out(par_done_reg249_out),
      .done(par_done_reg249_done)
  );
  
  std_reg #(1) par_done_reg250 (
      .in(par_done_reg250_in),
      .write_en(par_done_reg250_write_en),
      .clk(clk),
      .out(par_done_reg250_out),
      .done(par_done_reg250_done)
  );
  
  std_reg #(1) par_done_reg251 (
      .in(par_done_reg251_in),
      .write_en(par_done_reg251_write_en),
      .clk(clk),
      .out(par_done_reg251_out),
      .done(par_done_reg251_done)
  );
  
  std_reg #(1) par_done_reg252 (
      .in(par_done_reg252_in),
      .write_en(par_done_reg252_write_en),
      .clk(clk),
      .out(par_done_reg252_out),
      .done(par_done_reg252_done)
  );
  
  std_reg #(1) par_done_reg253 (
      .in(par_done_reg253_in),
      .write_en(par_done_reg253_write_en),
      .clk(clk),
      .out(par_done_reg253_out),
      .done(par_done_reg253_done)
  );
  
  std_reg #(1) par_done_reg254 (
      .in(par_done_reg254_in),
      .write_en(par_done_reg254_write_en),
      .clk(clk),
      .out(par_done_reg254_out),
      .done(par_done_reg254_done)
  );
  
  std_reg #(1) par_done_reg255 (
      .in(par_done_reg255_in),
      .write_en(par_done_reg255_write_en),
      .clk(clk),
      .out(par_done_reg255_out),
      .done(par_done_reg255_done)
  );
  
  std_reg #(1) par_done_reg256 (
      .in(par_done_reg256_in),
      .write_en(par_done_reg256_write_en),
      .clk(clk),
      .out(par_done_reg256_out),
      .done(par_done_reg256_done)
  );
  
  std_reg #(1) par_done_reg257 (
      .in(par_done_reg257_in),
      .write_en(par_done_reg257_write_en),
      .clk(clk),
      .out(par_done_reg257_out),
      .done(par_done_reg257_done)
  );
  
  std_reg #(1) par_done_reg258 (
      .in(par_done_reg258_in),
      .write_en(par_done_reg258_write_en),
      .clk(clk),
      .out(par_done_reg258_out),
      .done(par_done_reg258_done)
  );
  
  std_reg #(1) par_done_reg259 (
      .in(par_done_reg259_in),
      .write_en(par_done_reg259_write_en),
      .clk(clk),
      .out(par_done_reg259_out),
      .done(par_done_reg259_done)
  );
  
  std_reg #(1) par_done_reg260 (
      .in(par_done_reg260_in),
      .write_en(par_done_reg260_write_en),
      .clk(clk),
      .out(par_done_reg260_out),
      .done(par_done_reg260_done)
  );
  
  std_reg #(1) par_done_reg261 (
      .in(par_done_reg261_in),
      .write_en(par_done_reg261_write_en),
      .clk(clk),
      .out(par_done_reg261_out),
      .done(par_done_reg261_done)
  );
  
  std_reg #(1) par_done_reg262 (
      .in(par_done_reg262_in),
      .write_en(par_done_reg262_write_en),
      .clk(clk),
      .out(par_done_reg262_out),
      .done(par_done_reg262_done)
  );
  
  std_reg #(1) par_done_reg263 (
      .in(par_done_reg263_in),
      .write_en(par_done_reg263_write_en),
      .clk(clk),
      .out(par_done_reg263_out),
      .done(par_done_reg263_done)
  );
  
  std_reg #(1) par_done_reg264 (
      .in(par_done_reg264_in),
      .write_en(par_done_reg264_write_en),
      .clk(clk),
      .out(par_done_reg264_out),
      .done(par_done_reg264_done)
  );
  
  std_reg #(1) par_done_reg265 (
      .in(par_done_reg265_in),
      .write_en(par_done_reg265_write_en),
      .clk(clk),
      .out(par_done_reg265_out),
      .done(par_done_reg265_done)
  );
  
  std_reg #(1) par_done_reg266 (
      .in(par_done_reg266_in),
      .write_en(par_done_reg266_write_en),
      .clk(clk),
      .out(par_done_reg266_out),
      .done(par_done_reg266_done)
  );
  
  std_reg #(1) par_done_reg267 (
      .in(par_done_reg267_in),
      .write_en(par_done_reg267_write_en),
      .clk(clk),
      .out(par_done_reg267_out),
      .done(par_done_reg267_done)
  );
  
  std_reg #(1) par_done_reg268 (
      .in(par_done_reg268_in),
      .write_en(par_done_reg268_write_en),
      .clk(clk),
      .out(par_done_reg268_out),
      .done(par_done_reg268_done)
  );
  
  std_reg #(1) par_done_reg269 (
      .in(par_done_reg269_in),
      .write_en(par_done_reg269_write_en),
      .clk(clk),
      .out(par_done_reg269_out),
      .done(par_done_reg269_done)
  );
  
  std_reg #(1) par_done_reg270 (
      .in(par_done_reg270_in),
      .write_en(par_done_reg270_write_en),
      .clk(clk),
      .out(par_done_reg270_out),
      .done(par_done_reg270_done)
  );
  
  std_reg #(1) par_done_reg271 (
      .in(par_done_reg271_in),
      .write_en(par_done_reg271_write_en),
      .clk(clk),
      .out(par_done_reg271_out),
      .done(par_done_reg271_done)
  );
  
  std_reg #(1) par_done_reg272 (
      .in(par_done_reg272_in),
      .write_en(par_done_reg272_write_en),
      .clk(clk),
      .out(par_done_reg272_out),
      .done(par_done_reg272_done)
  );
  
  std_reg #(1) par_done_reg273 (
      .in(par_done_reg273_in),
      .write_en(par_done_reg273_write_en),
      .clk(clk),
      .out(par_done_reg273_out),
      .done(par_done_reg273_done)
  );
  
  std_reg #(1) par_done_reg274 (
      .in(par_done_reg274_in),
      .write_en(par_done_reg274_write_en),
      .clk(clk),
      .out(par_done_reg274_out),
      .done(par_done_reg274_done)
  );
  
  std_reg #(1) par_done_reg275 (
      .in(par_done_reg275_in),
      .write_en(par_done_reg275_write_en),
      .clk(clk),
      .out(par_done_reg275_out),
      .done(par_done_reg275_done)
  );
  
  std_reg #(1) par_done_reg276 (
      .in(par_done_reg276_in),
      .write_en(par_done_reg276_write_en),
      .clk(clk),
      .out(par_done_reg276_out),
      .done(par_done_reg276_done)
  );
  
  std_reg #(1) par_done_reg277 (
      .in(par_done_reg277_in),
      .write_en(par_done_reg277_write_en),
      .clk(clk),
      .out(par_done_reg277_out),
      .done(par_done_reg277_done)
  );
  
  std_reg #(1) par_done_reg278 (
      .in(par_done_reg278_in),
      .write_en(par_done_reg278_write_en),
      .clk(clk),
      .out(par_done_reg278_out),
      .done(par_done_reg278_done)
  );
  
  std_reg #(1) par_done_reg279 (
      .in(par_done_reg279_in),
      .write_en(par_done_reg279_write_en),
      .clk(clk),
      .out(par_done_reg279_out),
      .done(par_done_reg279_done)
  );
  
  std_reg #(1) par_done_reg280 (
      .in(par_done_reg280_in),
      .write_en(par_done_reg280_write_en),
      .clk(clk),
      .out(par_done_reg280_out),
      .done(par_done_reg280_done)
  );
  
  std_reg #(1) par_done_reg281 (
      .in(par_done_reg281_in),
      .write_en(par_done_reg281_write_en),
      .clk(clk),
      .out(par_done_reg281_out),
      .done(par_done_reg281_done)
  );
  
  std_reg #(1) par_done_reg282 (
      .in(par_done_reg282_in),
      .write_en(par_done_reg282_write_en),
      .clk(clk),
      .out(par_done_reg282_out),
      .done(par_done_reg282_done)
  );
  
  std_reg #(1) par_done_reg283 (
      .in(par_done_reg283_in),
      .write_en(par_done_reg283_write_en),
      .clk(clk),
      .out(par_done_reg283_out),
      .done(par_done_reg283_done)
  );
  
  std_reg #(1) par_done_reg284 (
      .in(par_done_reg284_in),
      .write_en(par_done_reg284_write_en),
      .clk(clk),
      .out(par_done_reg284_out),
      .done(par_done_reg284_done)
  );
  
  std_reg #(1) par_done_reg285 (
      .in(par_done_reg285_in),
      .write_en(par_done_reg285_write_en),
      .clk(clk),
      .out(par_done_reg285_out),
      .done(par_done_reg285_done)
  );
  
  std_reg #(1) par_done_reg286 (
      .in(par_done_reg286_in),
      .write_en(par_done_reg286_write_en),
      .clk(clk),
      .out(par_done_reg286_out),
      .done(par_done_reg286_done)
  );
  
  std_reg #(1) par_done_reg287 (
      .in(par_done_reg287_in),
      .write_en(par_done_reg287_write_en),
      .clk(clk),
      .out(par_done_reg287_out),
      .done(par_done_reg287_done)
  );
  
  std_reg #(1) par_done_reg288 (
      .in(par_done_reg288_in),
      .write_en(par_done_reg288_write_en),
      .clk(clk),
      .out(par_done_reg288_out),
      .done(par_done_reg288_done)
  );
  
  std_reg #(1) par_done_reg289 (
      .in(par_done_reg289_in),
      .write_en(par_done_reg289_write_en),
      .clk(clk),
      .out(par_done_reg289_out),
      .done(par_done_reg289_done)
  );
  
  std_reg #(1) par_done_reg290 (
      .in(par_done_reg290_in),
      .write_en(par_done_reg290_write_en),
      .clk(clk),
      .out(par_done_reg290_out),
      .done(par_done_reg290_done)
  );
  
  std_reg #(1) par_done_reg291 (
      .in(par_done_reg291_in),
      .write_en(par_done_reg291_write_en),
      .clk(clk),
      .out(par_done_reg291_out),
      .done(par_done_reg291_done)
  );
  
  std_reg #(1) par_done_reg292 (
      .in(par_done_reg292_in),
      .write_en(par_done_reg292_write_en),
      .clk(clk),
      .out(par_done_reg292_out),
      .done(par_done_reg292_done)
  );
  
  std_reg #(1) par_done_reg293 (
      .in(par_done_reg293_in),
      .write_en(par_done_reg293_write_en),
      .clk(clk),
      .out(par_done_reg293_out),
      .done(par_done_reg293_done)
  );
  
  std_reg #(1) par_done_reg294 (
      .in(par_done_reg294_in),
      .write_en(par_done_reg294_write_en),
      .clk(clk),
      .out(par_done_reg294_out),
      .done(par_done_reg294_done)
  );
  
  std_reg #(1) par_done_reg295 (
      .in(par_done_reg295_in),
      .write_en(par_done_reg295_write_en),
      .clk(clk),
      .out(par_done_reg295_out),
      .done(par_done_reg295_done)
  );
  
  std_reg #(1) par_reset15 (
      .in(par_reset15_in),
      .write_en(par_reset15_write_en),
      .clk(clk),
      .out(par_reset15_out),
      .done(par_reset15_done)
  );
  
  std_reg #(1) par_done_reg296 (
      .in(par_done_reg296_in),
      .write_en(par_done_reg296_write_en),
      .clk(clk),
      .out(par_done_reg296_out),
      .done(par_done_reg296_done)
  );
  
  std_reg #(1) par_done_reg297 (
      .in(par_done_reg297_in),
      .write_en(par_done_reg297_write_en),
      .clk(clk),
      .out(par_done_reg297_out),
      .done(par_done_reg297_done)
  );
  
  std_reg #(1) par_done_reg298 (
      .in(par_done_reg298_in),
      .write_en(par_done_reg298_write_en),
      .clk(clk),
      .out(par_done_reg298_out),
      .done(par_done_reg298_done)
  );
  
  std_reg #(1) par_done_reg299 (
      .in(par_done_reg299_in),
      .write_en(par_done_reg299_write_en),
      .clk(clk),
      .out(par_done_reg299_out),
      .done(par_done_reg299_done)
  );
  
  std_reg #(1) par_done_reg300 (
      .in(par_done_reg300_in),
      .write_en(par_done_reg300_write_en),
      .clk(clk),
      .out(par_done_reg300_out),
      .done(par_done_reg300_done)
  );
  
  std_reg #(1) par_done_reg301 (
      .in(par_done_reg301_in),
      .write_en(par_done_reg301_write_en),
      .clk(clk),
      .out(par_done_reg301_out),
      .done(par_done_reg301_done)
  );
  
  std_reg #(1) par_done_reg302 (
      .in(par_done_reg302_in),
      .write_en(par_done_reg302_write_en),
      .clk(clk),
      .out(par_done_reg302_out),
      .done(par_done_reg302_done)
  );
  
  std_reg #(1) par_done_reg303 (
      .in(par_done_reg303_in),
      .write_en(par_done_reg303_write_en),
      .clk(clk),
      .out(par_done_reg303_out),
      .done(par_done_reg303_done)
  );
  
  std_reg #(1) par_done_reg304 (
      .in(par_done_reg304_in),
      .write_en(par_done_reg304_write_en),
      .clk(clk),
      .out(par_done_reg304_out),
      .done(par_done_reg304_done)
  );
  
  std_reg #(1) par_done_reg305 (
      .in(par_done_reg305_in),
      .write_en(par_done_reg305_write_en),
      .clk(clk),
      .out(par_done_reg305_out),
      .done(par_done_reg305_done)
  );
  
  std_reg #(1) par_done_reg306 (
      .in(par_done_reg306_in),
      .write_en(par_done_reg306_write_en),
      .clk(clk),
      .out(par_done_reg306_out),
      .done(par_done_reg306_done)
  );
  
  std_reg #(1) par_done_reg307 (
      .in(par_done_reg307_in),
      .write_en(par_done_reg307_write_en),
      .clk(clk),
      .out(par_done_reg307_out),
      .done(par_done_reg307_done)
  );
  
  std_reg #(1) par_done_reg308 (
      .in(par_done_reg308_in),
      .write_en(par_done_reg308_write_en),
      .clk(clk),
      .out(par_done_reg308_out),
      .done(par_done_reg308_done)
  );
  
  std_reg #(1) par_done_reg309 (
      .in(par_done_reg309_in),
      .write_en(par_done_reg309_write_en),
      .clk(clk),
      .out(par_done_reg309_out),
      .done(par_done_reg309_done)
  );
  
  std_reg #(1) par_done_reg310 (
      .in(par_done_reg310_in),
      .write_en(par_done_reg310_write_en),
      .clk(clk),
      .out(par_done_reg310_out),
      .done(par_done_reg310_done)
  );
  
  std_reg #(1) par_done_reg311 (
      .in(par_done_reg311_in),
      .write_en(par_done_reg311_write_en),
      .clk(clk),
      .out(par_done_reg311_out),
      .done(par_done_reg311_done)
  );
  
  std_reg #(1) par_done_reg312 (
      .in(par_done_reg312_in),
      .write_en(par_done_reg312_write_en),
      .clk(clk),
      .out(par_done_reg312_out),
      .done(par_done_reg312_done)
  );
  
  std_reg #(1) par_done_reg313 (
      .in(par_done_reg313_in),
      .write_en(par_done_reg313_write_en),
      .clk(clk),
      .out(par_done_reg313_out),
      .done(par_done_reg313_done)
  );
  
  std_reg #(1) par_done_reg314 (
      .in(par_done_reg314_in),
      .write_en(par_done_reg314_write_en),
      .clk(clk),
      .out(par_done_reg314_out),
      .done(par_done_reg314_done)
  );
  
  std_reg #(1) par_done_reg315 (
      .in(par_done_reg315_in),
      .write_en(par_done_reg315_write_en),
      .clk(clk),
      .out(par_done_reg315_out),
      .done(par_done_reg315_done)
  );
  
  std_reg #(1) par_done_reg316 (
      .in(par_done_reg316_in),
      .write_en(par_done_reg316_write_en),
      .clk(clk),
      .out(par_done_reg316_out),
      .done(par_done_reg316_done)
  );
  
  std_reg #(1) par_done_reg317 (
      .in(par_done_reg317_in),
      .write_en(par_done_reg317_write_en),
      .clk(clk),
      .out(par_done_reg317_out),
      .done(par_done_reg317_done)
  );
  
  std_reg #(1) par_done_reg318 (
      .in(par_done_reg318_in),
      .write_en(par_done_reg318_write_en),
      .clk(clk),
      .out(par_done_reg318_out),
      .done(par_done_reg318_done)
  );
  
  std_reg #(1) par_done_reg319 (
      .in(par_done_reg319_in),
      .write_en(par_done_reg319_write_en),
      .clk(clk),
      .out(par_done_reg319_out),
      .done(par_done_reg319_done)
  );
  
  std_reg #(1) par_done_reg320 (
      .in(par_done_reg320_in),
      .write_en(par_done_reg320_write_en),
      .clk(clk),
      .out(par_done_reg320_out),
      .done(par_done_reg320_done)
  );
  
  std_reg #(1) par_done_reg321 (
      .in(par_done_reg321_in),
      .write_en(par_done_reg321_write_en),
      .clk(clk),
      .out(par_done_reg321_out),
      .done(par_done_reg321_done)
  );
  
  std_reg #(1) par_done_reg322 (
      .in(par_done_reg322_in),
      .write_en(par_done_reg322_write_en),
      .clk(clk),
      .out(par_done_reg322_out),
      .done(par_done_reg322_done)
  );
  
  std_reg #(1) par_done_reg323 (
      .in(par_done_reg323_in),
      .write_en(par_done_reg323_write_en),
      .clk(clk),
      .out(par_done_reg323_out),
      .done(par_done_reg323_done)
  );
  
  std_reg #(1) par_done_reg324 (
      .in(par_done_reg324_in),
      .write_en(par_done_reg324_write_en),
      .clk(clk),
      .out(par_done_reg324_out),
      .done(par_done_reg324_done)
  );
  
  std_reg #(1) par_done_reg325 (
      .in(par_done_reg325_in),
      .write_en(par_done_reg325_write_en),
      .clk(clk),
      .out(par_done_reg325_out),
      .done(par_done_reg325_done)
  );
  
  std_reg #(1) par_done_reg326 (
      .in(par_done_reg326_in),
      .write_en(par_done_reg326_write_en),
      .clk(clk),
      .out(par_done_reg326_out),
      .done(par_done_reg326_done)
  );
  
  std_reg #(1) par_done_reg327 (
      .in(par_done_reg327_in),
      .write_en(par_done_reg327_write_en),
      .clk(clk),
      .out(par_done_reg327_out),
      .done(par_done_reg327_done)
  );
  
  std_reg #(1) par_done_reg328 (
      .in(par_done_reg328_in),
      .write_en(par_done_reg328_write_en),
      .clk(clk),
      .out(par_done_reg328_out),
      .done(par_done_reg328_done)
  );
  
  std_reg #(1) par_done_reg329 (
      .in(par_done_reg329_in),
      .write_en(par_done_reg329_write_en),
      .clk(clk),
      .out(par_done_reg329_out),
      .done(par_done_reg329_done)
  );
  
  std_reg #(1) par_done_reg330 (
      .in(par_done_reg330_in),
      .write_en(par_done_reg330_write_en),
      .clk(clk),
      .out(par_done_reg330_out),
      .done(par_done_reg330_done)
  );
  
  std_reg #(1) par_done_reg331 (
      .in(par_done_reg331_in),
      .write_en(par_done_reg331_write_en),
      .clk(clk),
      .out(par_done_reg331_out),
      .done(par_done_reg331_done)
  );
  
  std_reg #(1) par_done_reg332 (
      .in(par_done_reg332_in),
      .write_en(par_done_reg332_write_en),
      .clk(clk),
      .out(par_done_reg332_out),
      .done(par_done_reg332_done)
  );
  
  std_reg #(1) par_done_reg333 (
      .in(par_done_reg333_in),
      .write_en(par_done_reg333_write_en),
      .clk(clk),
      .out(par_done_reg333_out),
      .done(par_done_reg333_done)
  );
  
  std_reg #(1) par_done_reg334 (
      .in(par_done_reg334_in),
      .write_en(par_done_reg334_write_en),
      .clk(clk),
      .out(par_done_reg334_out),
      .done(par_done_reg334_done)
  );
  
  std_reg #(1) par_done_reg335 (
      .in(par_done_reg335_in),
      .write_en(par_done_reg335_write_en),
      .clk(clk),
      .out(par_done_reg335_out),
      .done(par_done_reg335_done)
  );
  
  std_reg #(1) par_done_reg336 (
      .in(par_done_reg336_in),
      .write_en(par_done_reg336_write_en),
      .clk(clk),
      .out(par_done_reg336_out),
      .done(par_done_reg336_done)
  );
  
  std_reg #(1) par_done_reg337 (
      .in(par_done_reg337_in),
      .write_en(par_done_reg337_write_en),
      .clk(clk),
      .out(par_done_reg337_out),
      .done(par_done_reg337_done)
  );
  
  std_reg #(1) par_done_reg338 (
      .in(par_done_reg338_in),
      .write_en(par_done_reg338_write_en),
      .clk(clk),
      .out(par_done_reg338_out),
      .done(par_done_reg338_done)
  );
  
  std_reg #(1) par_done_reg339 (
      .in(par_done_reg339_in),
      .write_en(par_done_reg339_write_en),
      .clk(clk),
      .out(par_done_reg339_out),
      .done(par_done_reg339_done)
  );
  
  std_reg #(1) par_reset16 (
      .in(par_reset16_in),
      .write_en(par_reset16_write_en),
      .clk(clk),
      .out(par_reset16_out),
      .done(par_reset16_done)
  );
  
  std_reg #(1) par_done_reg340 (
      .in(par_done_reg340_in),
      .write_en(par_done_reg340_write_en),
      .clk(clk),
      .out(par_done_reg340_out),
      .done(par_done_reg340_done)
  );
  
  std_reg #(1) par_done_reg341 (
      .in(par_done_reg341_in),
      .write_en(par_done_reg341_write_en),
      .clk(clk),
      .out(par_done_reg341_out),
      .done(par_done_reg341_done)
  );
  
  std_reg #(1) par_done_reg342 (
      .in(par_done_reg342_in),
      .write_en(par_done_reg342_write_en),
      .clk(clk),
      .out(par_done_reg342_out),
      .done(par_done_reg342_done)
  );
  
  std_reg #(1) par_done_reg343 (
      .in(par_done_reg343_in),
      .write_en(par_done_reg343_write_en),
      .clk(clk),
      .out(par_done_reg343_out),
      .done(par_done_reg343_done)
  );
  
  std_reg #(1) par_done_reg344 (
      .in(par_done_reg344_in),
      .write_en(par_done_reg344_write_en),
      .clk(clk),
      .out(par_done_reg344_out),
      .done(par_done_reg344_done)
  );
  
  std_reg #(1) par_done_reg345 (
      .in(par_done_reg345_in),
      .write_en(par_done_reg345_write_en),
      .clk(clk),
      .out(par_done_reg345_out),
      .done(par_done_reg345_done)
  );
  
  std_reg #(1) par_done_reg346 (
      .in(par_done_reg346_in),
      .write_en(par_done_reg346_write_en),
      .clk(clk),
      .out(par_done_reg346_out),
      .done(par_done_reg346_done)
  );
  
  std_reg #(1) par_done_reg347 (
      .in(par_done_reg347_in),
      .write_en(par_done_reg347_write_en),
      .clk(clk),
      .out(par_done_reg347_out),
      .done(par_done_reg347_done)
  );
  
  std_reg #(1) par_done_reg348 (
      .in(par_done_reg348_in),
      .write_en(par_done_reg348_write_en),
      .clk(clk),
      .out(par_done_reg348_out),
      .done(par_done_reg348_done)
  );
  
  std_reg #(1) par_done_reg349 (
      .in(par_done_reg349_in),
      .write_en(par_done_reg349_write_en),
      .clk(clk),
      .out(par_done_reg349_out),
      .done(par_done_reg349_done)
  );
  
  std_reg #(1) par_done_reg350 (
      .in(par_done_reg350_in),
      .write_en(par_done_reg350_write_en),
      .clk(clk),
      .out(par_done_reg350_out),
      .done(par_done_reg350_done)
  );
  
  std_reg #(1) par_done_reg351 (
      .in(par_done_reg351_in),
      .write_en(par_done_reg351_write_en),
      .clk(clk),
      .out(par_done_reg351_out),
      .done(par_done_reg351_done)
  );
  
  std_reg #(1) par_done_reg352 (
      .in(par_done_reg352_in),
      .write_en(par_done_reg352_write_en),
      .clk(clk),
      .out(par_done_reg352_out),
      .done(par_done_reg352_done)
  );
  
  std_reg #(1) par_done_reg353 (
      .in(par_done_reg353_in),
      .write_en(par_done_reg353_write_en),
      .clk(clk),
      .out(par_done_reg353_out),
      .done(par_done_reg353_done)
  );
  
  std_reg #(1) par_done_reg354 (
      .in(par_done_reg354_in),
      .write_en(par_done_reg354_write_en),
      .clk(clk),
      .out(par_done_reg354_out),
      .done(par_done_reg354_done)
  );
  
  std_reg #(1) par_done_reg355 (
      .in(par_done_reg355_in),
      .write_en(par_done_reg355_write_en),
      .clk(clk),
      .out(par_done_reg355_out),
      .done(par_done_reg355_done)
  );
  
  std_reg #(1) par_done_reg356 (
      .in(par_done_reg356_in),
      .write_en(par_done_reg356_write_en),
      .clk(clk),
      .out(par_done_reg356_out),
      .done(par_done_reg356_done)
  );
  
  std_reg #(1) par_done_reg357 (
      .in(par_done_reg357_in),
      .write_en(par_done_reg357_write_en),
      .clk(clk),
      .out(par_done_reg357_out),
      .done(par_done_reg357_done)
  );
  
  std_reg #(1) par_done_reg358 (
      .in(par_done_reg358_in),
      .write_en(par_done_reg358_write_en),
      .clk(clk),
      .out(par_done_reg358_out),
      .done(par_done_reg358_done)
  );
  
  std_reg #(1) par_done_reg359 (
      .in(par_done_reg359_in),
      .write_en(par_done_reg359_write_en),
      .clk(clk),
      .out(par_done_reg359_out),
      .done(par_done_reg359_done)
  );
  
  std_reg #(1) par_done_reg360 (
      .in(par_done_reg360_in),
      .write_en(par_done_reg360_write_en),
      .clk(clk),
      .out(par_done_reg360_out),
      .done(par_done_reg360_done)
  );
  
  std_reg #(1) par_done_reg361 (
      .in(par_done_reg361_in),
      .write_en(par_done_reg361_write_en),
      .clk(clk),
      .out(par_done_reg361_out),
      .done(par_done_reg361_done)
  );
  
  std_reg #(1) par_done_reg362 (
      .in(par_done_reg362_in),
      .write_en(par_done_reg362_write_en),
      .clk(clk),
      .out(par_done_reg362_out),
      .done(par_done_reg362_done)
  );
  
  std_reg #(1) par_done_reg363 (
      .in(par_done_reg363_in),
      .write_en(par_done_reg363_write_en),
      .clk(clk),
      .out(par_done_reg363_out),
      .done(par_done_reg363_done)
  );
  
  std_reg #(1) par_done_reg364 (
      .in(par_done_reg364_in),
      .write_en(par_done_reg364_write_en),
      .clk(clk),
      .out(par_done_reg364_out),
      .done(par_done_reg364_done)
  );
  
  std_reg #(1) par_done_reg365 (
      .in(par_done_reg365_in),
      .write_en(par_done_reg365_write_en),
      .clk(clk),
      .out(par_done_reg365_out),
      .done(par_done_reg365_done)
  );
  
  std_reg #(1) par_done_reg366 (
      .in(par_done_reg366_in),
      .write_en(par_done_reg366_write_en),
      .clk(clk),
      .out(par_done_reg366_out),
      .done(par_done_reg366_done)
  );
  
  std_reg #(1) par_done_reg367 (
      .in(par_done_reg367_in),
      .write_en(par_done_reg367_write_en),
      .clk(clk),
      .out(par_done_reg367_out),
      .done(par_done_reg367_done)
  );
  
  std_reg #(1) par_done_reg368 (
      .in(par_done_reg368_in),
      .write_en(par_done_reg368_write_en),
      .clk(clk),
      .out(par_done_reg368_out),
      .done(par_done_reg368_done)
  );
  
  std_reg #(1) par_done_reg369 (
      .in(par_done_reg369_in),
      .write_en(par_done_reg369_write_en),
      .clk(clk),
      .out(par_done_reg369_out),
      .done(par_done_reg369_done)
  );
  
  std_reg #(1) par_done_reg370 (
      .in(par_done_reg370_in),
      .write_en(par_done_reg370_write_en),
      .clk(clk),
      .out(par_done_reg370_out),
      .done(par_done_reg370_done)
  );
  
  std_reg #(1) par_done_reg371 (
      .in(par_done_reg371_in),
      .write_en(par_done_reg371_write_en),
      .clk(clk),
      .out(par_done_reg371_out),
      .done(par_done_reg371_done)
  );
  
  std_reg #(1) par_done_reg372 (
      .in(par_done_reg372_in),
      .write_en(par_done_reg372_write_en),
      .clk(clk),
      .out(par_done_reg372_out),
      .done(par_done_reg372_done)
  );
  
  std_reg #(1) par_done_reg373 (
      .in(par_done_reg373_in),
      .write_en(par_done_reg373_write_en),
      .clk(clk),
      .out(par_done_reg373_out),
      .done(par_done_reg373_done)
  );
  
  std_reg #(1) par_done_reg374 (
      .in(par_done_reg374_in),
      .write_en(par_done_reg374_write_en),
      .clk(clk),
      .out(par_done_reg374_out),
      .done(par_done_reg374_done)
  );
  
  std_reg #(1) par_done_reg375 (
      .in(par_done_reg375_in),
      .write_en(par_done_reg375_write_en),
      .clk(clk),
      .out(par_done_reg375_out),
      .done(par_done_reg375_done)
  );
  
  std_reg #(1) par_done_reg376 (
      .in(par_done_reg376_in),
      .write_en(par_done_reg376_write_en),
      .clk(clk),
      .out(par_done_reg376_out),
      .done(par_done_reg376_done)
  );
  
  std_reg #(1) par_done_reg377 (
      .in(par_done_reg377_in),
      .write_en(par_done_reg377_write_en),
      .clk(clk),
      .out(par_done_reg377_out),
      .done(par_done_reg377_done)
  );
  
  std_reg #(1) par_done_reg378 (
      .in(par_done_reg378_in),
      .write_en(par_done_reg378_write_en),
      .clk(clk),
      .out(par_done_reg378_out),
      .done(par_done_reg378_done)
  );
  
  std_reg #(1) par_done_reg379 (
      .in(par_done_reg379_in),
      .write_en(par_done_reg379_write_en),
      .clk(clk),
      .out(par_done_reg379_out),
      .done(par_done_reg379_done)
  );
  
  std_reg #(1) par_done_reg380 (
      .in(par_done_reg380_in),
      .write_en(par_done_reg380_write_en),
      .clk(clk),
      .out(par_done_reg380_out),
      .done(par_done_reg380_done)
  );
  
  std_reg #(1) par_done_reg381 (
      .in(par_done_reg381_in),
      .write_en(par_done_reg381_write_en),
      .clk(clk),
      .out(par_done_reg381_out),
      .done(par_done_reg381_done)
  );
  
  std_reg #(1) par_done_reg382 (
      .in(par_done_reg382_in),
      .write_en(par_done_reg382_write_en),
      .clk(clk),
      .out(par_done_reg382_out),
      .done(par_done_reg382_done)
  );
  
  std_reg #(1) par_done_reg383 (
      .in(par_done_reg383_in),
      .write_en(par_done_reg383_write_en),
      .clk(clk),
      .out(par_done_reg383_out),
      .done(par_done_reg383_done)
  );
  
  std_reg #(1) par_done_reg384 (
      .in(par_done_reg384_in),
      .write_en(par_done_reg384_write_en),
      .clk(clk),
      .out(par_done_reg384_out),
      .done(par_done_reg384_done)
  );
  
  std_reg #(1) par_done_reg385 (
      .in(par_done_reg385_in),
      .write_en(par_done_reg385_write_en),
      .clk(clk),
      .out(par_done_reg385_out),
      .done(par_done_reg385_done)
  );
  
  std_reg #(1) par_done_reg386 (
      .in(par_done_reg386_in),
      .write_en(par_done_reg386_write_en),
      .clk(clk),
      .out(par_done_reg386_out),
      .done(par_done_reg386_done)
  );
  
  std_reg #(1) par_done_reg387 (
      .in(par_done_reg387_in),
      .write_en(par_done_reg387_write_en),
      .clk(clk),
      .out(par_done_reg387_out),
      .done(par_done_reg387_done)
  );
  
  std_reg #(1) par_done_reg388 (
      .in(par_done_reg388_in),
      .write_en(par_done_reg388_write_en),
      .clk(clk),
      .out(par_done_reg388_out),
      .done(par_done_reg388_done)
  );
  
  std_reg #(1) par_done_reg389 (
      .in(par_done_reg389_in),
      .write_en(par_done_reg389_write_en),
      .clk(clk),
      .out(par_done_reg389_out),
      .done(par_done_reg389_done)
  );
  
  std_reg #(1) par_done_reg390 (
      .in(par_done_reg390_in),
      .write_en(par_done_reg390_write_en),
      .clk(clk),
      .out(par_done_reg390_out),
      .done(par_done_reg390_done)
  );
  
  std_reg #(1) par_done_reg391 (
      .in(par_done_reg391_in),
      .write_en(par_done_reg391_write_en),
      .clk(clk),
      .out(par_done_reg391_out),
      .done(par_done_reg391_done)
  );
  
  std_reg #(1) par_done_reg392 (
      .in(par_done_reg392_in),
      .write_en(par_done_reg392_write_en),
      .clk(clk),
      .out(par_done_reg392_out),
      .done(par_done_reg392_done)
  );
  
  std_reg #(1) par_done_reg393 (
      .in(par_done_reg393_in),
      .write_en(par_done_reg393_write_en),
      .clk(clk),
      .out(par_done_reg393_out),
      .done(par_done_reg393_done)
  );
  
  std_reg #(1) par_done_reg394 (
      .in(par_done_reg394_in),
      .write_en(par_done_reg394_write_en),
      .clk(clk),
      .out(par_done_reg394_out),
      .done(par_done_reg394_done)
  );
  
  std_reg #(1) par_done_reg395 (
      .in(par_done_reg395_in),
      .write_en(par_done_reg395_write_en),
      .clk(clk),
      .out(par_done_reg395_out),
      .done(par_done_reg395_done)
  );
  
  std_reg #(1) par_done_reg396 (
      .in(par_done_reg396_in),
      .write_en(par_done_reg396_write_en),
      .clk(clk),
      .out(par_done_reg396_out),
      .done(par_done_reg396_done)
  );
  
  std_reg #(1) par_done_reg397 (
      .in(par_done_reg397_in),
      .write_en(par_done_reg397_write_en),
      .clk(clk),
      .out(par_done_reg397_out),
      .done(par_done_reg397_done)
  );
  
  std_reg #(1) par_done_reg398 (
      .in(par_done_reg398_in),
      .write_en(par_done_reg398_write_en),
      .clk(clk),
      .out(par_done_reg398_out),
      .done(par_done_reg398_done)
  );
  
  std_reg #(1) par_done_reg399 (
      .in(par_done_reg399_in),
      .write_en(par_done_reg399_write_en),
      .clk(clk),
      .out(par_done_reg399_out),
      .done(par_done_reg399_done)
  );
  
  std_reg #(1) par_done_reg400 (
      .in(par_done_reg400_in),
      .write_en(par_done_reg400_write_en),
      .clk(clk),
      .out(par_done_reg400_out),
      .done(par_done_reg400_done)
  );
  
  std_reg #(1) par_done_reg401 (
      .in(par_done_reg401_in),
      .write_en(par_done_reg401_write_en),
      .clk(clk),
      .out(par_done_reg401_out),
      .done(par_done_reg401_done)
  );
  
  std_reg #(1) par_done_reg402 (
      .in(par_done_reg402_in),
      .write_en(par_done_reg402_write_en),
      .clk(clk),
      .out(par_done_reg402_out),
      .done(par_done_reg402_done)
  );
  
  std_reg #(1) par_done_reg403 (
      .in(par_done_reg403_in),
      .write_en(par_done_reg403_write_en),
      .clk(clk),
      .out(par_done_reg403_out),
      .done(par_done_reg403_done)
  );
  
  std_reg #(1) par_done_reg404 (
      .in(par_done_reg404_in),
      .write_en(par_done_reg404_write_en),
      .clk(clk),
      .out(par_done_reg404_out),
      .done(par_done_reg404_done)
  );
  
  std_reg #(1) par_done_reg405 (
      .in(par_done_reg405_in),
      .write_en(par_done_reg405_write_en),
      .clk(clk),
      .out(par_done_reg405_out),
      .done(par_done_reg405_done)
  );
  
  std_reg #(1) par_done_reg406 (
      .in(par_done_reg406_in),
      .write_en(par_done_reg406_write_en),
      .clk(clk),
      .out(par_done_reg406_out),
      .done(par_done_reg406_done)
  );
  
  std_reg #(1) par_done_reg407 (
      .in(par_done_reg407_in),
      .write_en(par_done_reg407_write_en),
      .clk(clk),
      .out(par_done_reg407_out),
      .done(par_done_reg407_done)
  );
  
  std_reg #(1) par_done_reg408 (
      .in(par_done_reg408_in),
      .write_en(par_done_reg408_write_en),
      .clk(clk),
      .out(par_done_reg408_out),
      .done(par_done_reg408_done)
  );
  
  std_reg #(1) par_done_reg409 (
      .in(par_done_reg409_in),
      .write_en(par_done_reg409_write_en),
      .clk(clk),
      .out(par_done_reg409_out),
      .done(par_done_reg409_done)
  );
  
  std_reg #(1) par_done_reg410 (
      .in(par_done_reg410_in),
      .write_en(par_done_reg410_write_en),
      .clk(clk),
      .out(par_done_reg410_out),
      .done(par_done_reg410_done)
  );
  
  std_reg #(1) par_done_reg411 (
      .in(par_done_reg411_in),
      .write_en(par_done_reg411_write_en),
      .clk(clk),
      .out(par_done_reg411_out),
      .done(par_done_reg411_done)
  );
  
  std_reg #(1) par_reset17 (
      .in(par_reset17_in),
      .write_en(par_reset17_write_en),
      .clk(clk),
      .out(par_reset17_out),
      .done(par_reset17_done)
  );
  
  std_reg #(1) par_done_reg412 (
      .in(par_done_reg412_in),
      .write_en(par_done_reg412_write_en),
      .clk(clk),
      .out(par_done_reg412_out),
      .done(par_done_reg412_done)
  );
  
  std_reg #(1) par_done_reg413 (
      .in(par_done_reg413_in),
      .write_en(par_done_reg413_write_en),
      .clk(clk),
      .out(par_done_reg413_out),
      .done(par_done_reg413_done)
  );
  
  std_reg #(1) par_done_reg414 (
      .in(par_done_reg414_in),
      .write_en(par_done_reg414_write_en),
      .clk(clk),
      .out(par_done_reg414_out),
      .done(par_done_reg414_done)
  );
  
  std_reg #(1) par_done_reg415 (
      .in(par_done_reg415_in),
      .write_en(par_done_reg415_write_en),
      .clk(clk),
      .out(par_done_reg415_out),
      .done(par_done_reg415_done)
  );
  
  std_reg #(1) par_done_reg416 (
      .in(par_done_reg416_in),
      .write_en(par_done_reg416_write_en),
      .clk(clk),
      .out(par_done_reg416_out),
      .done(par_done_reg416_done)
  );
  
  std_reg #(1) par_done_reg417 (
      .in(par_done_reg417_in),
      .write_en(par_done_reg417_write_en),
      .clk(clk),
      .out(par_done_reg417_out),
      .done(par_done_reg417_done)
  );
  
  std_reg #(1) par_done_reg418 (
      .in(par_done_reg418_in),
      .write_en(par_done_reg418_write_en),
      .clk(clk),
      .out(par_done_reg418_out),
      .done(par_done_reg418_done)
  );
  
  std_reg #(1) par_done_reg419 (
      .in(par_done_reg419_in),
      .write_en(par_done_reg419_write_en),
      .clk(clk),
      .out(par_done_reg419_out),
      .done(par_done_reg419_done)
  );
  
  std_reg #(1) par_done_reg420 (
      .in(par_done_reg420_in),
      .write_en(par_done_reg420_write_en),
      .clk(clk),
      .out(par_done_reg420_out),
      .done(par_done_reg420_done)
  );
  
  std_reg #(1) par_done_reg421 (
      .in(par_done_reg421_in),
      .write_en(par_done_reg421_write_en),
      .clk(clk),
      .out(par_done_reg421_out),
      .done(par_done_reg421_done)
  );
  
  std_reg #(1) par_done_reg422 (
      .in(par_done_reg422_in),
      .write_en(par_done_reg422_write_en),
      .clk(clk),
      .out(par_done_reg422_out),
      .done(par_done_reg422_done)
  );
  
  std_reg #(1) par_done_reg423 (
      .in(par_done_reg423_in),
      .write_en(par_done_reg423_write_en),
      .clk(clk),
      .out(par_done_reg423_out),
      .done(par_done_reg423_done)
  );
  
  std_reg #(1) par_done_reg424 (
      .in(par_done_reg424_in),
      .write_en(par_done_reg424_write_en),
      .clk(clk),
      .out(par_done_reg424_out),
      .done(par_done_reg424_done)
  );
  
  std_reg #(1) par_done_reg425 (
      .in(par_done_reg425_in),
      .write_en(par_done_reg425_write_en),
      .clk(clk),
      .out(par_done_reg425_out),
      .done(par_done_reg425_done)
  );
  
  std_reg #(1) par_done_reg426 (
      .in(par_done_reg426_in),
      .write_en(par_done_reg426_write_en),
      .clk(clk),
      .out(par_done_reg426_out),
      .done(par_done_reg426_done)
  );
  
  std_reg #(1) par_done_reg427 (
      .in(par_done_reg427_in),
      .write_en(par_done_reg427_write_en),
      .clk(clk),
      .out(par_done_reg427_out),
      .done(par_done_reg427_done)
  );
  
  std_reg #(1) par_done_reg428 (
      .in(par_done_reg428_in),
      .write_en(par_done_reg428_write_en),
      .clk(clk),
      .out(par_done_reg428_out),
      .done(par_done_reg428_done)
  );
  
  std_reg #(1) par_done_reg429 (
      .in(par_done_reg429_in),
      .write_en(par_done_reg429_write_en),
      .clk(clk),
      .out(par_done_reg429_out),
      .done(par_done_reg429_done)
  );
  
  std_reg #(1) par_done_reg430 (
      .in(par_done_reg430_in),
      .write_en(par_done_reg430_write_en),
      .clk(clk),
      .out(par_done_reg430_out),
      .done(par_done_reg430_done)
  );
  
  std_reg #(1) par_done_reg431 (
      .in(par_done_reg431_in),
      .write_en(par_done_reg431_write_en),
      .clk(clk),
      .out(par_done_reg431_out),
      .done(par_done_reg431_done)
  );
  
  std_reg #(1) par_done_reg432 (
      .in(par_done_reg432_in),
      .write_en(par_done_reg432_write_en),
      .clk(clk),
      .out(par_done_reg432_out),
      .done(par_done_reg432_done)
  );
  
  std_reg #(1) par_done_reg433 (
      .in(par_done_reg433_in),
      .write_en(par_done_reg433_write_en),
      .clk(clk),
      .out(par_done_reg433_out),
      .done(par_done_reg433_done)
  );
  
  std_reg #(1) par_done_reg434 (
      .in(par_done_reg434_in),
      .write_en(par_done_reg434_write_en),
      .clk(clk),
      .out(par_done_reg434_out),
      .done(par_done_reg434_done)
  );
  
  std_reg #(1) par_done_reg435 (
      .in(par_done_reg435_in),
      .write_en(par_done_reg435_write_en),
      .clk(clk),
      .out(par_done_reg435_out),
      .done(par_done_reg435_done)
  );
  
  std_reg #(1) par_done_reg436 (
      .in(par_done_reg436_in),
      .write_en(par_done_reg436_write_en),
      .clk(clk),
      .out(par_done_reg436_out),
      .done(par_done_reg436_done)
  );
  
  std_reg #(1) par_done_reg437 (
      .in(par_done_reg437_in),
      .write_en(par_done_reg437_write_en),
      .clk(clk),
      .out(par_done_reg437_out),
      .done(par_done_reg437_done)
  );
  
  std_reg #(1) par_done_reg438 (
      .in(par_done_reg438_in),
      .write_en(par_done_reg438_write_en),
      .clk(clk),
      .out(par_done_reg438_out),
      .done(par_done_reg438_done)
  );
  
  std_reg #(1) par_done_reg439 (
      .in(par_done_reg439_in),
      .write_en(par_done_reg439_write_en),
      .clk(clk),
      .out(par_done_reg439_out),
      .done(par_done_reg439_done)
  );
  
  std_reg #(1) par_done_reg440 (
      .in(par_done_reg440_in),
      .write_en(par_done_reg440_write_en),
      .clk(clk),
      .out(par_done_reg440_out),
      .done(par_done_reg440_done)
  );
  
  std_reg #(1) par_done_reg441 (
      .in(par_done_reg441_in),
      .write_en(par_done_reg441_write_en),
      .clk(clk),
      .out(par_done_reg441_out),
      .done(par_done_reg441_done)
  );
  
  std_reg #(1) par_done_reg442 (
      .in(par_done_reg442_in),
      .write_en(par_done_reg442_write_en),
      .clk(clk),
      .out(par_done_reg442_out),
      .done(par_done_reg442_done)
  );
  
  std_reg #(1) par_done_reg443 (
      .in(par_done_reg443_in),
      .write_en(par_done_reg443_write_en),
      .clk(clk),
      .out(par_done_reg443_out),
      .done(par_done_reg443_done)
  );
  
  std_reg #(1) par_done_reg444 (
      .in(par_done_reg444_in),
      .write_en(par_done_reg444_write_en),
      .clk(clk),
      .out(par_done_reg444_out),
      .done(par_done_reg444_done)
  );
  
  std_reg #(1) par_done_reg445 (
      .in(par_done_reg445_in),
      .write_en(par_done_reg445_write_en),
      .clk(clk),
      .out(par_done_reg445_out),
      .done(par_done_reg445_done)
  );
  
  std_reg #(1) par_done_reg446 (
      .in(par_done_reg446_in),
      .write_en(par_done_reg446_write_en),
      .clk(clk),
      .out(par_done_reg446_out),
      .done(par_done_reg446_done)
  );
  
  std_reg #(1) par_done_reg447 (
      .in(par_done_reg447_in),
      .write_en(par_done_reg447_write_en),
      .clk(clk),
      .out(par_done_reg447_out),
      .done(par_done_reg447_done)
  );
  
  std_reg #(1) par_done_reg448 (
      .in(par_done_reg448_in),
      .write_en(par_done_reg448_write_en),
      .clk(clk),
      .out(par_done_reg448_out),
      .done(par_done_reg448_done)
  );
  
  std_reg #(1) par_done_reg449 (
      .in(par_done_reg449_in),
      .write_en(par_done_reg449_write_en),
      .clk(clk),
      .out(par_done_reg449_out),
      .done(par_done_reg449_done)
  );
  
  std_reg #(1) par_done_reg450 (
      .in(par_done_reg450_in),
      .write_en(par_done_reg450_write_en),
      .clk(clk),
      .out(par_done_reg450_out),
      .done(par_done_reg450_done)
  );
  
  std_reg #(1) par_done_reg451 (
      .in(par_done_reg451_in),
      .write_en(par_done_reg451_write_en),
      .clk(clk),
      .out(par_done_reg451_out),
      .done(par_done_reg451_done)
  );
  
  std_reg #(1) par_done_reg452 (
      .in(par_done_reg452_in),
      .write_en(par_done_reg452_write_en),
      .clk(clk),
      .out(par_done_reg452_out),
      .done(par_done_reg452_done)
  );
  
  std_reg #(1) par_done_reg453 (
      .in(par_done_reg453_in),
      .write_en(par_done_reg453_write_en),
      .clk(clk),
      .out(par_done_reg453_out),
      .done(par_done_reg453_done)
  );
  
  std_reg #(1) par_done_reg454 (
      .in(par_done_reg454_in),
      .write_en(par_done_reg454_write_en),
      .clk(clk),
      .out(par_done_reg454_out),
      .done(par_done_reg454_done)
  );
  
  std_reg #(1) par_done_reg455 (
      .in(par_done_reg455_in),
      .write_en(par_done_reg455_write_en),
      .clk(clk),
      .out(par_done_reg455_out),
      .done(par_done_reg455_done)
  );
  
  std_reg #(1) par_done_reg456 (
      .in(par_done_reg456_in),
      .write_en(par_done_reg456_write_en),
      .clk(clk),
      .out(par_done_reg456_out),
      .done(par_done_reg456_done)
  );
  
  std_reg #(1) par_done_reg457 (
      .in(par_done_reg457_in),
      .write_en(par_done_reg457_write_en),
      .clk(clk),
      .out(par_done_reg457_out),
      .done(par_done_reg457_done)
  );
  
  std_reg #(1) par_done_reg458 (
      .in(par_done_reg458_in),
      .write_en(par_done_reg458_write_en),
      .clk(clk),
      .out(par_done_reg458_out),
      .done(par_done_reg458_done)
  );
  
  std_reg #(1) par_done_reg459 (
      .in(par_done_reg459_in),
      .write_en(par_done_reg459_write_en),
      .clk(clk),
      .out(par_done_reg459_out),
      .done(par_done_reg459_done)
  );
  
  std_reg #(1) par_done_reg460 (
      .in(par_done_reg460_in),
      .write_en(par_done_reg460_write_en),
      .clk(clk),
      .out(par_done_reg460_out),
      .done(par_done_reg460_done)
  );
  
  std_reg #(1) par_done_reg461 (
      .in(par_done_reg461_in),
      .write_en(par_done_reg461_write_en),
      .clk(clk),
      .out(par_done_reg461_out),
      .done(par_done_reg461_done)
  );
  
  std_reg #(1) par_reset18 (
      .in(par_reset18_in),
      .write_en(par_reset18_write_en),
      .clk(clk),
      .out(par_reset18_out),
      .done(par_reset18_done)
  );
  
  std_reg #(1) par_done_reg462 (
      .in(par_done_reg462_in),
      .write_en(par_done_reg462_write_en),
      .clk(clk),
      .out(par_done_reg462_out),
      .done(par_done_reg462_done)
  );
  
  std_reg #(1) par_done_reg463 (
      .in(par_done_reg463_in),
      .write_en(par_done_reg463_write_en),
      .clk(clk),
      .out(par_done_reg463_out),
      .done(par_done_reg463_done)
  );
  
  std_reg #(1) par_done_reg464 (
      .in(par_done_reg464_in),
      .write_en(par_done_reg464_write_en),
      .clk(clk),
      .out(par_done_reg464_out),
      .done(par_done_reg464_done)
  );
  
  std_reg #(1) par_done_reg465 (
      .in(par_done_reg465_in),
      .write_en(par_done_reg465_write_en),
      .clk(clk),
      .out(par_done_reg465_out),
      .done(par_done_reg465_done)
  );
  
  std_reg #(1) par_done_reg466 (
      .in(par_done_reg466_in),
      .write_en(par_done_reg466_write_en),
      .clk(clk),
      .out(par_done_reg466_out),
      .done(par_done_reg466_done)
  );
  
  std_reg #(1) par_done_reg467 (
      .in(par_done_reg467_in),
      .write_en(par_done_reg467_write_en),
      .clk(clk),
      .out(par_done_reg467_out),
      .done(par_done_reg467_done)
  );
  
  std_reg #(1) par_done_reg468 (
      .in(par_done_reg468_in),
      .write_en(par_done_reg468_write_en),
      .clk(clk),
      .out(par_done_reg468_out),
      .done(par_done_reg468_done)
  );
  
  std_reg #(1) par_done_reg469 (
      .in(par_done_reg469_in),
      .write_en(par_done_reg469_write_en),
      .clk(clk),
      .out(par_done_reg469_out),
      .done(par_done_reg469_done)
  );
  
  std_reg #(1) par_done_reg470 (
      .in(par_done_reg470_in),
      .write_en(par_done_reg470_write_en),
      .clk(clk),
      .out(par_done_reg470_out),
      .done(par_done_reg470_done)
  );
  
  std_reg #(1) par_done_reg471 (
      .in(par_done_reg471_in),
      .write_en(par_done_reg471_write_en),
      .clk(clk),
      .out(par_done_reg471_out),
      .done(par_done_reg471_done)
  );
  
  std_reg #(1) par_done_reg472 (
      .in(par_done_reg472_in),
      .write_en(par_done_reg472_write_en),
      .clk(clk),
      .out(par_done_reg472_out),
      .done(par_done_reg472_done)
  );
  
  std_reg #(1) par_done_reg473 (
      .in(par_done_reg473_in),
      .write_en(par_done_reg473_write_en),
      .clk(clk),
      .out(par_done_reg473_out),
      .done(par_done_reg473_done)
  );
  
  std_reg #(1) par_done_reg474 (
      .in(par_done_reg474_in),
      .write_en(par_done_reg474_write_en),
      .clk(clk),
      .out(par_done_reg474_out),
      .done(par_done_reg474_done)
  );
  
  std_reg #(1) par_done_reg475 (
      .in(par_done_reg475_in),
      .write_en(par_done_reg475_write_en),
      .clk(clk),
      .out(par_done_reg475_out),
      .done(par_done_reg475_done)
  );
  
  std_reg #(1) par_done_reg476 (
      .in(par_done_reg476_in),
      .write_en(par_done_reg476_write_en),
      .clk(clk),
      .out(par_done_reg476_out),
      .done(par_done_reg476_done)
  );
  
  std_reg #(1) par_done_reg477 (
      .in(par_done_reg477_in),
      .write_en(par_done_reg477_write_en),
      .clk(clk),
      .out(par_done_reg477_out),
      .done(par_done_reg477_done)
  );
  
  std_reg #(1) par_done_reg478 (
      .in(par_done_reg478_in),
      .write_en(par_done_reg478_write_en),
      .clk(clk),
      .out(par_done_reg478_out),
      .done(par_done_reg478_done)
  );
  
  std_reg #(1) par_done_reg479 (
      .in(par_done_reg479_in),
      .write_en(par_done_reg479_write_en),
      .clk(clk),
      .out(par_done_reg479_out),
      .done(par_done_reg479_done)
  );
  
  std_reg #(1) par_done_reg480 (
      .in(par_done_reg480_in),
      .write_en(par_done_reg480_write_en),
      .clk(clk),
      .out(par_done_reg480_out),
      .done(par_done_reg480_done)
  );
  
  std_reg #(1) par_done_reg481 (
      .in(par_done_reg481_in),
      .write_en(par_done_reg481_write_en),
      .clk(clk),
      .out(par_done_reg481_out),
      .done(par_done_reg481_done)
  );
  
  std_reg #(1) par_done_reg482 (
      .in(par_done_reg482_in),
      .write_en(par_done_reg482_write_en),
      .clk(clk),
      .out(par_done_reg482_out),
      .done(par_done_reg482_done)
  );
  
  std_reg #(1) par_done_reg483 (
      .in(par_done_reg483_in),
      .write_en(par_done_reg483_write_en),
      .clk(clk),
      .out(par_done_reg483_out),
      .done(par_done_reg483_done)
  );
  
  std_reg #(1) par_done_reg484 (
      .in(par_done_reg484_in),
      .write_en(par_done_reg484_write_en),
      .clk(clk),
      .out(par_done_reg484_out),
      .done(par_done_reg484_done)
  );
  
  std_reg #(1) par_done_reg485 (
      .in(par_done_reg485_in),
      .write_en(par_done_reg485_write_en),
      .clk(clk),
      .out(par_done_reg485_out),
      .done(par_done_reg485_done)
  );
  
  std_reg #(1) par_done_reg486 (
      .in(par_done_reg486_in),
      .write_en(par_done_reg486_write_en),
      .clk(clk),
      .out(par_done_reg486_out),
      .done(par_done_reg486_done)
  );
  
  std_reg #(1) par_done_reg487 (
      .in(par_done_reg487_in),
      .write_en(par_done_reg487_write_en),
      .clk(clk),
      .out(par_done_reg487_out),
      .done(par_done_reg487_done)
  );
  
  std_reg #(1) par_done_reg488 (
      .in(par_done_reg488_in),
      .write_en(par_done_reg488_write_en),
      .clk(clk),
      .out(par_done_reg488_out),
      .done(par_done_reg488_done)
  );
  
  std_reg #(1) par_done_reg489 (
      .in(par_done_reg489_in),
      .write_en(par_done_reg489_write_en),
      .clk(clk),
      .out(par_done_reg489_out),
      .done(par_done_reg489_done)
  );
  
  std_reg #(1) par_done_reg490 (
      .in(par_done_reg490_in),
      .write_en(par_done_reg490_write_en),
      .clk(clk),
      .out(par_done_reg490_out),
      .done(par_done_reg490_done)
  );
  
  std_reg #(1) par_done_reg491 (
      .in(par_done_reg491_in),
      .write_en(par_done_reg491_write_en),
      .clk(clk),
      .out(par_done_reg491_out),
      .done(par_done_reg491_done)
  );
  
  std_reg #(1) par_done_reg492 (
      .in(par_done_reg492_in),
      .write_en(par_done_reg492_write_en),
      .clk(clk),
      .out(par_done_reg492_out),
      .done(par_done_reg492_done)
  );
  
  std_reg #(1) par_done_reg493 (
      .in(par_done_reg493_in),
      .write_en(par_done_reg493_write_en),
      .clk(clk),
      .out(par_done_reg493_out),
      .done(par_done_reg493_done)
  );
  
  std_reg #(1) par_done_reg494 (
      .in(par_done_reg494_in),
      .write_en(par_done_reg494_write_en),
      .clk(clk),
      .out(par_done_reg494_out),
      .done(par_done_reg494_done)
  );
  
  std_reg #(1) par_done_reg495 (
      .in(par_done_reg495_in),
      .write_en(par_done_reg495_write_en),
      .clk(clk),
      .out(par_done_reg495_out),
      .done(par_done_reg495_done)
  );
  
  std_reg #(1) par_done_reg496 (
      .in(par_done_reg496_in),
      .write_en(par_done_reg496_write_en),
      .clk(clk),
      .out(par_done_reg496_out),
      .done(par_done_reg496_done)
  );
  
  std_reg #(1) par_done_reg497 (
      .in(par_done_reg497_in),
      .write_en(par_done_reg497_write_en),
      .clk(clk),
      .out(par_done_reg497_out),
      .done(par_done_reg497_done)
  );
  
  std_reg #(1) par_done_reg498 (
      .in(par_done_reg498_in),
      .write_en(par_done_reg498_write_en),
      .clk(clk),
      .out(par_done_reg498_out),
      .done(par_done_reg498_done)
  );
  
  std_reg #(1) par_done_reg499 (
      .in(par_done_reg499_in),
      .write_en(par_done_reg499_write_en),
      .clk(clk),
      .out(par_done_reg499_out),
      .done(par_done_reg499_done)
  );
  
  std_reg #(1) par_done_reg500 (
      .in(par_done_reg500_in),
      .write_en(par_done_reg500_write_en),
      .clk(clk),
      .out(par_done_reg500_out),
      .done(par_done_reg500_done)
  );
  
  std_reg #(1) par_done_reg501 (
      .in(par_done_reg501_in),
      .write_en(par_done_reg501_write_en),
      .clk(clk),
      .out(par_done_reg501_out),
      .done(par_done_reg501_done)
  );
  
  std_reg #(1) par_done_reg502 (
      .in(par_done_reg502_in),
      .write_en(par_done_reg502_write_en),
      .clk(clk),
      .out(par_done_reg502_out),
      .done(par_done_reg502_done)
  );
  
  std_reg #(1) par_done_reg503 (
      .in(par_done_reg503_in),
      .write_en(par_done_reg503_write_en),
      .clk(clk),
      .out(par_done_reg503_out),
      .done(par_done_reg503_done)
  );
  
  std_reg #(1) par_done_reg504 (
      .in(par_done_reg504_in),
      .write_en(par_done_reg504_write_en),
      .clk(clk),
      .out(par_done_reg504_out),
      .done(par_done_reg504_done)
  );
  
  std_reg #(1) par_done_reg505 (
      .in(par_done_reg505_in),
      .write_en(par_done_reg505_write_en),
      .clk(clk),
      .out(par_done_reg505_out),
      .done(par_done_reg505_done)
  );
  
  std_reg #(1) par_done_reg506 (
      .in(par_done_reg506_in),
      .write_en(par_done_reg506_write_en),
      .clk(clk),
      .out(par_done_reg506_out),
      .done(par_done_reg506_done)
  );
  
  std_reg #(1) par_done_reg507 (
      .in(par_done_reg507_in),
      .write_en(par_done_reg507_write_en),
      .clk(clk),
      .out(par_done_reg507_out),
      .done(par_done_reg507_done)
  );
  
  std_reg #(1) par_done_reg508 (
      .in(par_done_reg508_in),
      .write_en(par_done_reg508_write_en),
      .clk(clk),
      .out(par_done_reg508_out),
      .done(par_done_reg508_done)
  );
  
  std_reg #(1) par_done_reg509 (
      .in(par_done_reg509_in),
      .write_en(par_done_reg509_write_en),
      .clk(clk),
      .out(par_done_reg509_out),
      .done(par_done_reg509_done)
  );
  
  std_reg #(1) par_done_reg510 (
      .in(par_done_reg510_in),
      .write_en(par_done_reg510_write_en),
      .clk(clk),
      .out(par_done_reg510_out),
      .done(par_done_reg510_done)
  );
  
  std_reg #(1) par_done_reg511 (
      .in(par_done_reg511_in),
      .write_en(par_done_reg511_write_en),
      .clk(clk),
      .out(par_done_reg511_out),
      .done(par_done_reg511_done)
  );
  
  std_reg #(1) par_done_reg512 (
      .in(par_done_reg512_in),
      .write_en(par_done_reg512_write_en),
      .clk(clk),
      .out(par_done_reg512_out),
      .done(par_done_reg512_done)
  );
  
  std_reg #(1) par_done_reg513 (
      .in(par_done_reg513_in),
      .write_en(par_done_reg513_write_en),
      .clk(clk),
      .out(par_done_reg513_out),
      .done(par_done_reg513_done)
  );
  
  std_reg #(1) par_done_reg514 (
      .in(par_done_reg514_in),
      .write_en(par_done_reg514_write_en),
      .clk(clk),
      .out(par_done_reg514_out),
      .done(par_done_reg514_done)
  );
  
  std_reg #(1) par_done_reg515 (
      .in(par_done_reg515_in),
      .write_en(par_done_reg515_write_en),
      .clk(clk),
      .out(par_done_reg515_out),
      .done(par_done_reg515_done)
  );
  
  std_reg #(1) par_done_reg516 (
      .in(par_done_reg516_in),
      .write_en(par_done_reg516_write_en),
      .clk(clk),
      .out(par_done_reg516_out),
      .done(par_done_reg516_done)
  );
  
  std_reg #(1) par_done_reg517 (
      .in(par_done_reg517_in),
      .write_en(par_done_reg517_write_en),
      .clk(clk),
      .out(par_done_reg517_out),
      .done(par_done_reg517_done)
  );
  
  std_reg #(1) par_done_reg518 (
      .in(par_done_reg518_in),
      .write_en(par_done_reg518_write_en),
      .clk(clk),
      .out(par_done_reg518_out),
      .done(par_done_reg518_done)
  );
  
  std_reg #(1) par_done_reg519 (
      .in(par_done_reg519_in),
      .write_en(par_done_reg519_write_en),
      .clk(clk),
      .out(par_done_reg519_out),
      .done(par_done_reg519_done)
  );
  
  std_reg #(1) par_done_reg520 (
      .in(par_done_reg520_in),
      .write_en(par_done_reg520_write_en),
      .clk(clk),
      .out(par_done_reg520_out),
      .done(par_done_reg520_done)
  );
  
  std_reg #(1) par_done_reg521 (
      .in(par_done_reg521_in),
      .write_en(par_done_reg521_write_en),
      .clk(clk),
      .out(par_done_reg521_out),
      .done(par_done_reg521_done)
  );
  
  std_reg #(1) par_done_reg522 (
      .in(par_done_reg522_in),
      .write_en(par_done_reg522_write_en),
      .clk(clk),
      .out(par_done_reg522_out),
      .done(par_done_reg522_done)
  );
  
  std_reg #(1) par_done_reg523 (
      .in(par_done_reg523_in),
      .write_en(par_done_reg523_write_en),
      .clk(clk),
      .out(par_done_reg523_out),
      .done(par_done_reg523_done)
  );
  
  std_reg #(1) par_done_reg524 (
      .in(par_done_reg524_in),
      .write_en(par_done_reg524_write_en),
      .clk(clk),
      .out(par_done_reg524_out),
      .done(par_done_reg524_done)
  );
  
  std_reg #(1) par_done_reg525 (
      .in(par_done_reg525_in),
      .write_en(par_done_reg525_write_en),
      .clk(clk),
      .out(par_done_reg525_out),
      .done(par_done_reg525_done)
  );
  
  std_reg #(1) par_done_reg526 (
      .in(par_done_reg526_in),
      .write_en(par_done_reg526_write_en),
      .clk(clk),
      .out(par_done_reg526_out),
      .done(par_done_reg526_done)
  );
  
  std_reg #(1) par_done_reg527 (
      .in(par_done_reg527_in),
      .write_en(par_done_reg527_write_en),
      .clk(clk),
      .out(par_done_reg527_out),
      .done(par_done_reg527_done)
  );
  
  std_reg #(1) par_done_reg528 (
      .in(par_done_reg528_in),
      .write_en(par_done_reg528_write_en),
      .clk(clk),
      .out(par_done_reg528_out),
      .done(par_done_reg528_done)
  );
  
  std_reg #(1) par_done_reg529 (
      .in(par_done_reg529_in),
      .write_en(par_done_reg529_write_en),
      .clk(clk),
      .out(par_done_reg529_out),
      .done(par_done_reg529_done)
  );
  
  std_reg #(1) par_done_reg530 (
      .in(par_done_reg530_in),
      .write_en(par_done_reg530_write_en),
      .clk(clk),
      .out(par_done_reg530_out),
      .done(par_done_reg530_done)
  );
  
  std_reg #(1) par_done_reg531 (
      .in(par_done_reg531_in),
      .write_en(par_done_reg531_write_en),
      .clk(clk),
      .out(par_done_reg531_out),
      .done(par_done_reg531_done)
  );
  
  std_reg #(1) par_done_reg532 (
      .in(par_done_reg532_in),
      .write_en(par_done_reg532_write_en),
      .clk(clk),
      .out(par_done_reg532_out),
      .done(par_done_reg532_done)
  );
  
  std_reg #(1) par_done_reg533 (
      .in(par_done_reg533_in),
      .write_en(par_done_reg533_write_en),
      .clk(clk),
      .out(par_done_reg533_out),
      .done(par_done_reg533_done)
  );
  
  std_reg #(1) par_done_reg534 (
      .in(par_done_reg534_in),
      .write_en(par_done_reg534_write_en),
      .clk(clk),
      .out(par_done_reg534_out),
      .done(par_done_reg534_done)
  );
  
  std_reg #(1) par_done_reg535 (
      .in(par_done_reg535_in),
      .write_en(par_done_reg535_write_en),
      .clk(clk),
      .out(par_done_reg535_out),
      .done(par_done_reg535_done)
  );
  
  std_reg #(1) par_done_reg536 (
      .in(par_done_reg536_in),
      .write_en(par_done_reg536_write_en),
      .clk(clk),
      .out(par_done_reg536_out),
      .done(par_done_reg536_done)
  );
  
  std_reg #(1) par_done_reg537 (
      .in(par_done_reg537_in),
      .write_en(par_done_reg537_write_en),
      .clk(clk),
      .out(par_done_reg537_out),
      .done(par_done_reg537_done)
  );
  
  std_reg #(1) par_done_reg538 (
      .in(par_done_reg538_in),
      .write_en(par_done_reg538_write_en),
      .clk(clk),
      .out(par_done_reg538_out),
      .done(par_done_reg538_done)
  );
  
  std_reg #(1) par_done_reg539 (
      .in(par_done_reg539_in),
      .write_en(par_done_reg539_write_en),
      .clk(clk),
      .out(par_done_reg539_out),
      .done(par_done_reg539_done)
  );
  
  std_reg #(1) par_done_reg540 (
      .in(par_done_reg540_in),
      .write_en(par_done_reg540_write_en),
      .clk(clk),
      .out(par_done_reg540_out),
      .done(par_done_reg540_done)
  );
  
  std_reg #(1) par_done_reg541 (
      .in(par_done_reg541_in),
      .write_en(par_done_reg541_write_en),
      .clk(clk),
      .out(par_done_reg541_out),
      .done(par_done_reg541_done)
  );
  
  std_reg #(1) par_done_reg542 (
      .in(par_done_reg542_in),
      .write_en(par_done_reg542_write_en),
      .clk(clk),
      .out(par_done_reg542_out),
      .done(par_done_reg542_done)
  );
  
  std_reg #(1) par_done_reg543 (
      .in(par_done_reg543_in),
      .write_en(par_done_reg543_write_en),
      .clk(clk),
      .out(par_done_reg543_out),
      .done(par_done_reg543_done)
  );
  
  std_reg #(1) par_done_reg544 (
      .in(par_done_reg544_in),
      .write_en(par_done_reg544_write_en),
      .clk(clk),
      .out(par_done_reg544_out),
      .done(par_done_reg544_done)
  );
  
  std_reg #(1) par_done_reg545 (
      .in(par_done_reg545_in),
      .write_en(par_done_reg545_write_en),
      .clk(clk),
      .out(par_done_reg545_out),
      .done(par_done_reg545_done)
  );
  
  std_reg #(1) par_reset19 (
      .in(par_reset19_in),
      .write_en(par_reset19_write_en),
      .clk(clk),
      .out(par_reset19_out),
      .done(par_reset19_done)
  );
  
  std_reg #(1) par_done_reg546 (
      .in(par_done_reg546_in),
      .write_en(par_done_reg546_write_en),
      .clk(clk),
      .out(par_done_reg546_out),
      .done(par_done_reg546_done)
  );
  
  std_reg #(1) par_done_reg547 (
      .in(par_done_reg547_in),
      .write_en(par_done_reg547_write_en),
      .clk(clk),
      .out(par_done_reg547_out),
      .done(par_done_reg547_done)
  );
  
  std_reg #(1) par_done_reg548 (
      .in(par_done_reg548_in),
      .write_en(par_done_reg548_write_en),
      .clk(clk),
      .out(par_done_reg548_out),
      .done(par_done_reg548_done)
  );
  
  std_reg #(1) par_done_reg549 (
      .in(par_done_reg549_in),
      .write_en(par_done_reg549_write_en),
      .clk(clk),
      .out(par_done_reg549_out),
      .done(par_done_reg549_done)
  );
  
  std_reg #(1) par_done_reg550 (
      .in(par_done_reg550_in),
      .write_en(par_done_reg550_write_en),
      .clk(clk),
      .out(par_done_reg550_out),
      .done(par_done_reg550_done)
  );
  
  std_reg #(1) par_done_reg551 (
      .in(par_done_reg551_in),
      .write_en(par_done_reg551_write_en),
      .clk(clk),
      .out(par_done_reg551_out),
      .done(par_done_reg551_done)
  );
  
  std_reg #(1) par_done_reg552 (
      .in(par_done_reg552_in),
      .write_en(par_done_reg552_write_en),
      .clk(clk),
      .out(par_done_reg552_out),
      .done(par_done_reg552_done)
  );
  
  std_reg #(1) par_done_reg553 (
      .in(par_done_reg553_in),
      .write_en(par_done_reg553_write_en),
      .clk(clk),
      .out(par_done_reg553_out),
      .done(par_done_reg553_done)
  );
  
  std_reg #(1) par_done_reg554 (
      .in(par_done_reg554_in),
      .write_en(par_done_reg554_write_en),
      .clk(clk),
      .out(par_done_reg554_out),
      .done(par_done_reg554_done)
  );
  
  std_reg #(1) par_done_reg555 (
      .in(par_done_reg555_in),
      .write_en(par_done_reg555_write_en),
      .clk(clk),
      .out(par_done_reg555_out),
      .done(par_done_reg555_done)
  );
  
  std_reg #(1) par_done_reg556 (
      .in(par_done_reg556_in),
      .write_en(par_done_reg556_write_en),
      .clk(clk),
      .out(par_done_reg556_out),
      .done(par_done_reg556_done)
  );
  
  std_reg #(1) par_done_reg557 (
      .in(par_done_reg557_in),
      .write_en(par_done_reg557_write_en),
      .clk(clk),
      .out(par_done_reg557_out),
      .done(par_done_reg557_done)
  );
  
  std_reg #(1) par_done_reg558 (
      .in(par_done_reg558_in),
      .write_en(par_done_reg558_write_en),
      .clk(clk),
      .out(par_done_reg558_out),
      .done(par_done_reg558_done)
  );
  
  std_reg #(1) par_done_reg559 (
      .in(par_done_reg559_in),
      .write_en(par_done_reg559_write_en),
      .clk(clk),
      .out(par_done_reg559_out),
      .done(par_done_reg559_done)
  );
  
  std_reg #(1) par_done_reg560 (
      .in(par_done_reg560_in),
      .write_en(par_done_reg560_write_en),
      .clk(clk),
      .out(par_done_reg560_out),
      .done(par_done_reg560_done)
  );
  
  std_reg #(1) par_done_reg561 (
      .in(par_done_reg561_in),
      .write_en(par_done_reg561_write_en),
      .clk(clk),
      .out(par_done_reg561_out),
      .done(par_done_reg561_done)
  );
  
  std_reg #(1) par_done_reg562 (
      .in(par_done_reg562_in),
      .write_en(par_done_reg562_write_en),
      .clk(clk),
      .out(par_done_reg562_out),
      .done(par_done_reg562_done)
  );
  
  std_reg #(1) par_done_reg563 (
      .in(par_done_reg563_in),
      .write_en(par_done_reg563_write_en),
      .clk(clk),
      .out(par_done_reg563_out),
      .done(par_done_reg563_done)
  );
  
  std_reg #(1) par_done_reg564 (
      .in(par_done_reg564_in),
      .write_en(par_done_reg564_write_en),
      .clk(clk),
      .out(par_done_reg564_out),
      .done(par_done_reg564_done)
  );
  
  std_reg #(1) par_done_reg565 (
      .in(par_done_reg565_in),
      .write_en(par_done_reg565_write_en),
      .clk(clk),
      .out(par_done_reg565_out),
      .done(par_done_reg565_done)
  );
  
  std_reg #(1) par_done_reg566 (
      .in(par_done_reg566_in),
      .write_en(par_done_reg566_write_en),
      .clk(clk),
      .out(par_done_reg566_out),
      .done(par_done_reg566_done)
  );
  
  std_reg #(1) par_done_reg567 (
      .in(par_done_reg567_in),
      .write_en(par_done_reg567_write_en),
      .clk(clk),
      .out(par_done_reg567_out),
      .done(par_done_reg567_done)
  );
  
  std_reg #(1) par_done_reg568 (
      .in(par_done_reg568_in),
      .write_en(par_done_reg568_write_en),
      .clk(clk),
      .out(par_done_reg568_out),
      .done(par_done_reg568_done)
  );
  
  std_reg #(1) par_done_reg569 (
      .in(par_done_reg569_in),
      .write_en(par_done_reg569_write_en),
      .clk(clk),
      .out(par_done_reg569_out),
      .done(par_done_reg569_done)
  );
  
  std_reg #(1) par_done_reg570 (
      .in(par_done_reg570_in),
      .write_en(par_done_reg570_write_en),
      .clk(clk),
      .out(par_done_reg570_out),
      .done(par_done_reg570_done)
  );
  
  std_reg #(1) par_done_reg571 (
      .in(par_done_reg571_in),
      .write_en(par_done_reg571_write_en),
      .clk(clk),
      .out(par_done_reg571_out),
      .done(par_done_reg571_done)
  );
  
  std_reg #(1) par_done_reg572 (
      .in(par_done_reg572_in),
      .write_en(par_done_reg572_write_en),
      .clk(clk),
      .out(par_done_reg572_out),
      .done(par_done_reg572_done)
  );
  
  std_reg #(1) par_done_reg573 (
      .in(par_done_reg573_in),
      .write_en(par_done_reg573_write_en),
      .clk(clk),
      .out(par_done_reg573_out),
      .done(par_done_reg573_done)
  );
  
  std_reg #(1) par_done_reg574 (
      .in(par_done_reg574_in),
      .write_en(par_done_reg574_write_en),
      .clk(clk),
      .out(par_done_reg574_out),
      .done(par_done_reg574_done)
  );
  
  std_reg #(1) par_done_reg575 (
      .in(par_done_reg575_in),
      .write_en(par_done_reg575_write_en),
      .clk(clk),
      .out(par_done_reg575_out),
      .done(par_done_reg575_done)
  );
  
  std_reg #(1) par_done_reg576 (
      .in(par_done_reg576_in),
      .write_en(par_done_reg576_write_en),
      .clk(clk),
      .out(par_done_reg576_out),
      .done(par_done_reg576_done)
  );
  
  std_reg #(1) par_done_reg577 (
      .in(par_done_reg577_in),
      .write_en(par_done_reg577_write_en),
      .clk(clk),
      .out(par_done_reg577_out),
      .done(par_done_reg577_done)
  );
  
  std_reg #(1) par_done_reg578 (
      .in(par_done_reg578_in),
      .write_en(par_done_reg578_write_en),
      .clk(clk),
      .out(par_done_reg578_out),
      .done(par_done_reg578_done)
  );
  
  std_reg #(1) par_done_reg579 (
      .in(par_done_reg579_in),
      .write_en(par_done_reg579_write_en),
      .clk(clk),
      .out(par_done_reg579_out),
      .done(par_done_reg579_done)
  );
  
  std_reg #(1) par_done_reg580 (
      .in(par_done_reg580_in),
      .write_en(par_done_reg580_write_en),
      .clk(clk),
      .out(par_done_reg580_out),
      .done(par_done_reg580_done)
  );
  
  std_reg #(1) par_done_reg581 (
      .in(par_done_reg581_in),
      .write_en(par_done_reg581_write_en),
      .clk(clk),
      .out(par_done_reg581_out),
      .done(par_done_reg581_done)
  );
  
  std_reg #(1) par_done_reg582 (
      .in(par_done_reg582_in),
      .write_en(par_done_reg582_write_en),
      .clk(clk),
      .out(par_done_reg582_out),
      .done(par_done_reg582_done)
  );
  
  std_reg #(1) par_done_reg583 (
      .in(par_done_reg583_in),
      .write_en(par_done_reg583_write_en),
      .clk(clk),
      .out(par_done_reg583_out),
      .done(par_done_reg583_done)
  );
  
  std_reg #(1) par_done_reg584 (
      .in(par_done_reg584_in),
      .write_en(par_done_reg584_write_en),
      .clk(clk),
      .out(par_done_reg584_out),
      .done(par_done_reg584_done)
  );
  
  std_reg #(1) par_done_reg585 (
      .in(par_done_reg585_in),
      .write_en(par_done_reg585_write_en),
      .clk(clk),
      .out(par_done_reg585_out),
      .done(par_done_reg585_done)
  );
  
  std_reg #(1) par_done_reg586 (
      .in(par_done_reg586_in),
      .write_en(par_done_reg586_write_en),
      .clk(clk),
      .out(par_done_reg586_out),
      .done(par_done_reg586_done)
  );
  
  std_reg #(1) par_done_reg587 (
      .in(par_done_reg587_in),
      .write_en(par_done_reg587_write_en),
      .clk(clk),
      .out(par_done_reg587_out),
      .done(par_done_reg587_done)
  );
  
  std_reg #(1) par_done_reg588 (
      .in(par_done_reg588_in),
      .write_en(par_done_reg588_write_en),
      .clk(clk),
      .out(par_done_reg588_out),
      .done(par_done_reg588_done)
  );
  
  std_reg #(1) par_done_reg589 (
      .in(par_done_reg589_in),
      .write_en(par_done_reg589_write_en),
      .clk(clk),
      .out(par_done_reg589_out),
      .done(par_done_reg589_done)
  );
  
  std_reg #(1) par_done_reg590 (
      .in(par_done_reg590_in),
      .write_en(par_done_reg590_write_en),
      .clk(clk),
      .out(par_done_reg590_out),
      .done(par_done_reg590_done)
  );
  
  std_reg #(1) par_done_reg591 (
      .in(par_done_reg591_in),
      .write_en(par_done_reg591_write_en),
      .clk(clk),
      .out(par_done_reg591_out),
      .done(par_done_reg591_done)
  );
  
  std_reg #(1) par_done_reg592 (
      .in(par_done_reg592_in),
      .write_en(par_done_reg592_write_en),
      .clk(clk),
      .out(par_done_reg592_out),
      .done(par_done_reg592_done)
  );
  
  std_reg #(1) par_done_reg593 (
      .in(par_done_reg593_in),
      .write_en(par_done_reg593_write_en),
      .clk(clk),
      .out(par_done_reg593_out),
      .done(par_done_reg593_done)
  );
  
  std_reg #(1) par_done_reg594 (
      .in(par_done_reg594_in),
      .write_en(par_done_reg594_write_en),
      .clk(clk),
      .out(par_done_reg594_out),
      .done(par_done_reg594_done)
  );
  
  std_reg #(1) par_done_reg595 (
      .in(par_done_reg595_in),
      .write_en(par_done_reg595_write_en),
      .clk(clk),
      .out(par_done_reg595_out),
      .done(par_done_reg595_done)
  );
  
  std_reg #(1) par_done_reg596 (
      .in(par_done_reg596_in),
      .write_en(par_done_reg596_write_en),
      .clk(clk),
      .out(par_done_reg596_out),
      .done(par_done_reg596_done)
  );
  
  std_reg #(1) par_done_reg597 (
      .in(par_done_reg597_in),
      .write_en(par_done_reg597_write_en),
      .clk(clk),
      .out(par_done_reg597_out),
      .done(par_done_reg597_done)
  );
  
  std_reg #(1) par_done_reg598 (
      .in(par_done_reg598_in),
      .write_en(par_done_reg598_write_en),
      .clk(clk),
      .out(par_done_reg598_out),
      .done(par_done_reg598_done)
  );
  
  std_reg #(1) par_done_reg599 (
      .in(par_done_reg599_in),
      .write_en(par_done_reg599_write_en),
      .clk(clk),
      .out(par_done_reg599_out),
      .done(par_done_reg599_done)
  );
  
  std_reg #(1) par_reset20 (
      .in(par_reset20_in),
      .write_en(par_reset20_write_en),
      .clk(clk),
      .out(par_reset20_out),
      .done(par_reset20_done)
  );
  
  std_reg #(1) par_done_reg600 (
      .in(par_done_reg600_in),
      .write_en(par_done_reg600_write_en),
      .clk(clk),
      .out(par_done_reg600_out),
      .done(par_done_reg600_done)
  );
  
  std_reg #(1) par_done_reg601 (
      .in(par_done_reg601_in),
      .write_en(par_done_reg601_write_en),
      .clk(clk),
      .out(par_done_reg601_out),
      .done(par_done_reg601_done)
  );
  
  std_reg #(1) par_done_reg602 (
      .in(par_done_reg602_in),
      .write_en(par_done_reg602_write_en),
      .clk(clk),
      .out(par_done_reg602_out),
      .done(par_done_reg602_done)
  );
  
  std_reg #(1) par_done_reg603 (
      .in(par_done_reg603_in),
      .write_en(par_done_reg603_write_en),
      .clk(clk),
      .out(par_done_reg603_out),
      .done(par_done_reg603_done)
  );
  
  std_reg #(1) par_done_reg604 (
      .in(par_done_reg604_in),
      .write_en(par_done_reg604_write_en),
      .clk(clk),
      .out(par_done_reg604_out),
      .done(par_done_reg604_done)
  );
  
  std_reg #(1) par_done_reg605 (
      .in(par_done_reg605_in),
      .write_en(par_done_reg605_write_en),
      .clk(clk),
      .out(par_done_reg605_out),
      .done(par_done_reg605_done)
  );
  
  std_reg #(1) par_done_reg606 (
      .in(par_done_reg606_in),
      .write_en(par_done_reg606_write_en),
      .clk(clk),
      .out(par_done_reg606_out),
      .done(par_done_reg606_done)
  );
  
  std_reg #(1) par_done_reg607 (
      .in(par_done_reg607_in),
      .write_en(par_done_reg607_write_en),
      .clk(clk),
      .out(par_done_reg607_out),
      .done(par_done_reg607_done)
  );
  
  std_reg #(1) par_done_reg608 (
      .in(par_done_reg608_in),
      .write_en(par_done_reg608_write_en),
      .clk(clk),
      .out(par_done_reg608_out),
      .done(par_done_reg608_done)
  );
  
  std_reg #(1) par_done_reg609 (
      .in(par_done_reg609_in),
      .write_en(par_done_reg609_write_en),
      .clk(clk),
      .out(par_done_reg609_out),
      .done(par_done_reg609_done)
  );
  
  std_reg #(1) par_done_reg610 (
      .in(par_done_reg610_in),
      .write_en(par_done_reg610_write_en),
      .clk(clk),
      .out(par_done_reg610_out),
      .done(par_done_reg610_done)
  );
  
  std_reg #(1) par_done_reg611 (
      .in(par_done_reg611_in),
      .write_en(par_done_reg611_write_en),
      .clk(clk),
      .out(par_done_reg611_out),
      .done(par_done_reg611_done)
  );
  
  std_reg #(1) par_done_reg612 (
      .in(par_done_reg612_in),
      .write_en(par_done_reg612_write_en),
      .clk(clk),
      .out(par_done_reg612_out),
      .done(par_done_reg612_done)
  );
  
  std_reg #(1) par_done_reg613 (
      .in(par_done_reg613_in),
      .write_en(par_done_reg613_write_en),
      .clk(clk),
      .out(par_done_reg613_out),
      .done(par_done_reg613_done)
  );
  
  std_reg #(1) par_done_reg614 (
      .in(par_done_reg614_in),
      .write_en(par_done_reg614_write_en),
      .clk(clk),
      .out(par_done_reg614_out),
      .done(par_done_reg614_done)
  );
  
  std_reg #(1) par_done_reg615 (
      .in(par_done_reg615_in),
      .write_en(par_done_reg615_write_en),
      .clk(clk),
      .out(par_done_reg615_out),
      .done(par_done_reg615_done)
  );
  
  std_reg #(1) par_done_reg616 (
      .in(par_done_reg616_in),
      .write_en(par_done_reg616_write_en),
      .clk(clk),
      .out(par_done_reg616_out),
      .done(par_done_reg616_done)
  );
  
  std_reg #(1) par_done_reg617 (
      .in(par_done_reg617_in),
      .write_en(par_done_reg617_write_en),
      .clk(clk),
      .out(par_done_reg617_out),
      .done(par_done_reg617_done)
  );
  
  std_reg #(1) par_done_reg618 (
      .in(par_done_reg618_in),
      .write_en(par_done_reg618_write_en),
      .clk(clk),
      .out(par_done_reg618_out),
      .done(par_done_reg618_done)
  );
  
  std_reg #(1) par_done_reg619 (
      .in(par_done_reg619_in),
      .write_en(par_done_reg619_write_en),
      .clk(clk),
      .out(par_done_reg619_out),
      .done(par_done_reg619_done)
  );
  
  std_reg #(1) par_done_reg620 (
      .in(par_done_reg620_in),
      .write_en(par_done_reg620_write_en),
      .clk(clk),
      .out(par_done_reg620_out),
      .done(par_done_reg620_done)
  );
  
  std_reg #(1) par_done_reg621 (
      .in(par_done_reg621_in),
      .write_en(par_done_reg621_write_en),
      .clk(clk),
      .out(par_done_reg621_out),
      .done(par_done_reg621_done)
  );
  
  std_reg #(1) par_done_reg622 (
      .in(par_done_reg622_in),
      .write_en(par_done_reg622_write_en),
      .clk(clk),
      .out(par_done_reg622_out),
      .done(par_done_reg622_done)
  );
  
  std_reg #(1) par_done_reg623 (
      .in(par_done_reg623_in),
      .write_en(par_done_reg623_write_en),
      .clk(clk),
      .out(par_done_reg623_out),
      .done(par_done_reg623_done)
  );
  
  std_reg #(1) par_done_reg624 (
      .in(par_done_reg624_in),
      .write_en(par_done_reg624_write_en),
      .clk(clk),
      .out(par_done_reg624_out),
      .done(par_done_reg624_done)
  );
  
  std_reg #(1) par_done_reg625 (
      .in(par_done_reg625_in),
      .write_en(par_done_reg625_write_en),
      .clk(clk),
      .out(par_done_reg625_out),
      .done(par_done_reg625_done)
  );
  
  std_reg #(1) par_done_reg626 (
      .in(par_done_reg626_in),
      .write_en(par_done_reg626_write_en),
      .clk(clk),
      .out(par_done_reg626_out),
      .done(par_done_reg626_done)
  );
  
  std_reg #(1) par_done_reg627 (
      .in(par_done_reg627_in),
      .write_en(par_done_reg627_write_en),
      .clk(clk),
      .out(par_done_reg627_out),
      .done(par_done_reg627_done)
  );
  
  std_reg #(1) par_done_reg628 (
      .in(par_done_reg628_in),
      .write_en(par_done_reg628_write_en),
      .clk(clk),
      .out(par_done_reg628_out),
      .done(par_done_reg628_done)
  );
  
  std_reg #(1) par_done_reg629 (
      .in(par_done_reg629_in),
      .write_en(par_done_reg629_write_en),
      .clk(clk),
      .out(par_done_reg629_out),
      .done(par_done_reg629_done)
  );
  
  std_reg #(1) par_done_reg630 (
      .in(par_done_reg630_in),
      .write_en(par_done_reg630_write_en),
      .clk(clk),
      .out(par_done_reg630_out),
      .done(par_done_reg630_done)
  );
  
  std_reg #(1) par_done_reg631 (
      .in(par_done_reg631_in),
      .write_en(par_done_reg631_write_en),
      .clk(clk),
      .out(par_done_reg631_out),
      .done(par_done_reg631_done)
  );
  
  std_reg #(1) par_done_reg632 (
      .in(par_done_reg632_in),
      .write_en(par_done_reg632_write_en),
      .clk(clk),
      .out(par_done_reg632_out),
      .done(par_done_reg632_done)
  );
  
  std_reg #(1) par_done_reg633 (
      .in(par_done_reg633_in),
      .write_en(par_done_reg633_write_en),
      .clk(clk),
      .out(par_done_reg633_out),
      .done(par_done_reg633_done)
  );
  
  std_reg #(1) par_done_reg634 (
      .in(par_done_reg634_in),
      .write_en(par_done_reg634_write_en),
      .clk(clk),
      .out(par_done_reg634_out),
      .done(par_done_reg634_done)
  );
  
  std_reg #(1) par_done_reg635 (
      .in(par_done_reg635_in),
      .write_en(par_done_reg635_write_en),
      .clk(clk),
      .out(par_done_reg635_out),
      .done(par_done_reg635_done)
  );
  
  std_reg #(1) par_done_reg636 (
      .in(par_done_reg636_in),
      .write_en(par_done_reg636_write_en),
      .clk(clk),
      .out(par_done_reg636_out),
      .done(par_done_reg636_done)
  );
  
  std_reg #(1) par_done_reg637 (
      .in(par_done_reg637_in),
      .write_en(par_done_reg637_write_en),
      .clk(clk),
      .out(par_done_reg637_out),
      .done(par_done_reg637_done)
  );
  
  std_reg #(1) par_done_reg638 (
      .in(par_done_reg638_in),
      .write_en(par_done_reg638_write_en),
      .clk(clk),
      .out(par_done_reg638_out),
      .done(par_done_reg638_done)
  );
  
  std_reg #(1) par_done_reg639 (
      .in(par_done_reg639_in),
      .write_en(par_done_reg639_write_en),
      .clk(clk),
      .out(par_done_reg639_out),
      .done(par_done_reg639_done)
  );
  
  std_reg #(1) par_done_reg640 (
      .in(par_done_reg640_in),
      .write_en(par_done_reg640_write_en),
      .clk(clk),
      .out(par_done_reg640_out),
      .done(par_done_reg640_done)
  );
  
  std_reg #(1) par_done_reg641 (
      .in(par_done_reg641_in),
      .write_en(par_done_reg641_write_en),
      .clk(clk),
      .out(par_done_reg641_out),
      .done(par_done_reg641_done)
  );
  
  std_reg #(1) par_done_reg642 (
      .in(par_done_reg642_in),
      .write_en(par_done_reg642_write_en),
      .clk(clk),
      .out(par_done_reg642_out),
      .done(par_done_reg642_done)
  );
  
  std_reg #(1) par_done_reg643 (
      .in(par_done_reg643_in),
      .write_en(par_done_reg643_write_en),
      .clk(clk),
      .out(par_done_reg643_out),
      .done(par_done_reg643_done)
  );
  
  std_reg #(1) par_done_reg644 (
      .in(par_done_reg644_in),
      .write_en(par_done_reg644_write_en),
      .clk(clk),
      .out(par_done_reg644_out),
      .done(par_done_reg644_done)
  );
  
  std_reg #(1) par_done_reg645 (
      .in(par_done_reg645_in),
      .write_en(par_done_reg645_write_en),
      .clk(clk),
      .out(par_done_reg645_out),
      .done(par_done_reg645_done)
  );
  
  std_reg #(1) par_done_reg646 (
      .in(par_done_reg646_in),
      .write_en(par_done_reg646_write_en),
      .clk(clk),
      .out(par_done_reg646_out),
      .done(par_done_reg646_done)
  );
  
  std_reg #(1) par_done_reg647 (
      .in(par_done_reg647_in),
      .write_en(par_done_reg647_write_en),
      .clk(clk),
      .out(par_done_reg647_out),
      .done(par_done_reg647_done)
  );
  
  std_reg #(1) par_done_reg648 (
      .in(par_done_reg648_in),
      .write_en(par_done_reg648_write_en),
      .clk(clk),
      .out(par_done_reg648_out),
      .done(par_done_reg648_done)
  );
  
  std_reg #(1) par_done_reg649 (
      .in(par_done_reg649_in),
      .write_en(par_done_reg649_write_en),
      .clk(clk),
      .out(par_done_reg649_out),
      .done(par_done_reg649_done)
  );
  
  std_reg #(1) par_done_reg650 (
      .in(par_done_reg650_in),
      .write_en(par_done_reg650_write_en),
      .clk(clk),
      .out(par_done_reg650_out),
      .done(par_done_reg650_done)
  );
  
  std_reg #(1) par_done_reg651 (
      .in(par_done_reg651_in),
      .write_en(par_done_reg651_write_en),
      .clk(clk),
      .out(par_done_reg651_out),
      .done(par_done_reg651_done)
  );
  
  std_reg #(1) par_done_reg652 (
      .in(par_done_reg652_in),
      .write_en(par_done_reg652_write_en),
      .clk(clk),
      .out(par_done_reg652_out),
      .done(par_done_reg652_done)
  );
  
  std_reg #(1) par_done_reg653 (
      .in(par_done_reg653_in),
      .write_en(par_done_reg653_write_en),
      .clk(clk),
      .out(par_done_reg653_out),
      .done(par_done_reg653_done)
  );
  
  std_reg #(1) par_done_reg654 (
      .in(par_done_reg654_in),
      .write_en(par_done_reg654_write_en),
      .clk(clk),
      .out(par_done_reg654_out),
      .done(par_done_reg654_done)
  );
  
  std_reg #(1) par_done_reg655 (
      .in(par_done_reg655_in),
      .write_en(par_done_reg655_write_en),
      .clk(clk),
      .out(par_done_reg655_out),
      .done(par_done_reg655_done)
  );
  
  std_reg #(1) par_done_reg656 (
      .in(par_done_reg656_in),
      .write_en(par_done_reg656_write_en),
      .clk(clk),
      .out(par_done_reg656_out),
      .done(par_done_reg656_done)
  );
  
  std_reg #(1) par_done_reg657 (
      .in(par_done_reg657_in),
      .write_en(par_done_reg657_write_en),
      .clk(clk),
      .out(par_done_reg657_out),
      .done(par_done_reg657_done)
  );
  
  std_reg #(1) par_done_reg658 (
      .in(par_done_reg658_in),
      .write_en(par_done_reg658_write_en),
      .clk(clk),
      .out(par_done_reg658_out),
      .done(par_done_reg658_done)
  );
  
  std_reg #(1) par_done_reg659 (
      .in(par_done_reg659_in),
      .write_en(par_done_reg659_write_en),
      .clk(clk),
      .out(par_done_reg659_out),
      .done(par_done_reg659_done)
  );
  
  std_reg #(1) par_done_reg660 (
      .in(par_done_reg660_in),
      .write_en(par_done_reg660_write_en),
      .clk(clk),
      .out(par_done_reg660_out),
      .done(par_done_reg660_done)
  );
  
  std_reg #(1) par_done_reg661 (
      .in(par_done_reg661_in),
      .write_en(par_done_reg661_write_en),
      .clk(clk),
      .out(par_done_reg661_out),
      .done(par_done_reg661_done)
  );
  
  std_reg #(1) par_done_reg662 (
      .in(par_done_reg662_in),
      .write_en(par_done_reg662_write_en),
      .clk(clk),
      .out(par_done_reg662_out),
      .done(par_done_reg662_done)
  );
  
  std_reg #(1) par_done_reg663 (
      .in(par_done_reg663_in),
      .write_en(par_done_reg663_write_en),
      .clk(clk),
      .out(par_done_reg663_out),
      .done(par_done_reg663_done)
  );
  
  std_reg #(1) par_done_reg664 (
      .in(par_done_reg664_in),
      .write_en(par_done_reg664_write_en),
      .clk(clk),
      .out(par_done_reg664_out),
      .done(par_done_reg664_done)
  );
  
  std_reg #(1) par_done_reg665 (
      .in(par_done_reg665_in),
      .write_en(par_done_reg665_write_en),
      .clk(clk),
      .out(par_done_reg665_out),
      .done(par_done_reg665_done)
  );
  
  std_reg #(1) par_done_reg666 (
      .in(par_done_reg666_in),
      .write_en(par_done_reg666_write_en),
      .clk(clk),
      .out(par_done_reg666_out),
      .done(par_done_reg666_done)
  );
  
  std_reg #(1) par_done_reg667 (
      .in(par_done_reg667_in),
      .write_en(par_done_reg667_write_en),
      .clk(clk),
      .out(par_done_reg667_out),
      .done(par_done_reg667_done)
  );
  
  std_reg #(1) par_done_reg668 (
      .in(par_done_reg668_in),
      .write_en(par_done_reg668_write_en),
      .clk(clk),
      .out(par_done_reg668_out),
      .done(par_done_reg668_done)
  );
  
  std_reg #(1) par_done_reg669 (
      .in(par_done_reg669_in),
      .write_en(par_done_reg669_write_en),
      .clk(clk),
      .out(par_done_reg669_out),
      .done(par_done_reg669_done)
  );
  
  std_reg #(1) par_done_reg670 (
      .in(par_done_reg670_in),
      .write_en(par_done_reg670_write_en),
      .clk(clk),
      .out(par_done_reg670_out),
      .done(par_done_reg670_done)
  );
  
  std_reg #(1) par_done_reg671 (
      .in(par_done_reg671_in),
      .write_en(par_done_reg671_write_en),
      .clk(clk),
      .out(par_done_reg671_out),
      .done(par_done_reg671_done)
  );
  
  std_reg #(1) par_done_reg672 (
      .in(par_done_reg672_in),
      .write_en(par_done_reg672_write_en),
      .clk(clk),
      .out(par_done_reg672_out),
      .done(par_done_reg672_done)
  );
  
  std_reg #(1) par_done_reg673 (
      .in(par_done_reg673_in),
      .write_en(par_done_reg673_write_en),
      .clk(clk),
      .out(par_done_reg673_out),
      .done(par_done_reg673_done)
  );
  
  std_reg #(1) par_done_reg674 (
      .in(par_done_reg674_in),
      .write_en(par_done_reg674_write_en),
      .clk(clk),
      .out(par_done_reg674_out),
      .done(par_done_reg674_done)
  );
  
  std_reg #(1) par_done_reg675 (
      .in(par_done_reg675_in),
      .write_en(par_done_reg675_write_en),
      .clk(clk),
      .out(par_done_reg675_out),
      .done(par_done_reg675_done)
  );
  
  std_reg #(1) par_done_reg676 (
      .in(par_done_reg676_in),
      .write_en(par_done_reg676_write_en),
      .clk(clk),
      .out(par_done_reg676_out),
      .done(par_done_reg676_done)
  );
  
  std_reg #(1) par_done_reg677 (
      .in(par_done_reg677_in),
      .write_en(par_done_reg677_write_en),
      .clk(clk),
      .out(par_done_reg677_out),
      .done(par_done_reg677_done)
  );
  
  std_reg #(1) par_done_reg678 (
      .in(par_done_reg678_in),
      .write_en(par_done_reg678_write_en),
      .clk(clk),
      .out(par_done_reg678_out),
      .done(par_done_reg678_done)
  );
  
  std_reg #(1) par_done_reg679 (
      .in(par_done_reg679_in),
      .write_en(par_done_reg679_write_en),
      .clk(clk),
      .out(par_done_reg679_out),
      .done(par_done_reg679_done)
  );
  
  std_reg #(1) par_done_reg680 (
      .in(par_done_reg680_in),
      .write_en(par_done_reg680_write_en),
      .clk(clk),
      .out(par_done_reg680_out),
      .done(par_done_reg680_done)
  );
  
  std_reg #(1) par_done_reg681 (
      .in(par_done_reg681_in),
      .write_en(par_done_reg681_write_en),
      .clk(clk),
      .out(par_done_reg681_out),
      .done(par_done_reg681_done)
  );
  
  std_reg #(1) par_done_reg682 (
      .in(par_done_reg682_in),
      .write_en(par_done_reg682_write_en),
      .clk(clk),
      .out(par_done_reg682_out),
      .done(par_done_reg682_done)
  );
  
  std_reg #(1) par_done_reg683 (
      .in(par_done_reg683_in),
      .write_en(par_done_reg683_write_en),
      .clk(clk),
      .out(par_done_reg683_out),
      .done(par_done_reg683_done)
  );
  
  std_reg #(1) par_done_reg684 (
      .in(par_done_reg684_in),
      .write_en(par_done_reg684_write_en),
      .clk(clk),
      .out(par_done_reg684_out),
      .done(par_done_reg684_done)
  );
  
  std_reg #(1) par_done_reg685 (
      .in(par_done_reg685_in),
      .write_en(par_done_reg685_write_en),
      .clk(clk),
      .out(par_done_reg685_out),
      .done(par_done_reg685_done)
  );
  
  std_reg #(1) par_done_reg686 (
      .in(par_done_reg686_in),
      .write_en(par_done_reg686_write_en),
      .clk(clk),
      .out(par_done_reg686_out),
      .done(par_done_reg686_done)
  );
  
  std_reg #(1) par_done_reg687 (
      .in(par_done_reg687_in),
      .write_en(par_done_reg687_write_en),
      .clk(clk),
      .out(par_done_reg687_out),
      .done(par_done_reg687_done)
  );
  
  std_reg #(1) par_done_reg688 (
      .in(par_done_reg688_in),
      .write_en(par_done_reg688_write_en),
      .clk(clk),
      .out(par_done_reg688_out),
      .done(par_done_reg688_done)
  );
  
  std_reg #(1) par_done_reg689 (
      .in(par_done_reg689_in),
      .write_en(par_done_reg689_write_en),
      .clk(clk),
      .out(par_done_reg689_out),
      .done(par_done_reg689_done)
  );
  
  std_reg #(1) par_done_reg690 (
      .in(par_done_reg690_in),
      .write_en(par_done_reg690_write_en),
      .clk(clk),
      .out(par_done_reg690_out),
      .done(par_done_reg690_done)
  );
  
  std_reg #(1) par_done_reg691 (
      .in(par_done_reg691_in),
      .write_en(par_done_reg691_write_en),
      .clk(clk),
      .out(par_done_reg691_out),
      .done(par_done_reg691_done)
  );
  
  std_reg #(1) par_reset21 (
      .in(par_reset21_in),
      .write_en(par_reset21_write_en),
      .clk(clk),
      .out(par_reset21_out),
      .done(par_reset21_done)
  );
  
  std_reg #(1) par_done_reg692 (
      .in(par_done_reg692_in),
      .write_en(par_done_reg692_write_en),
      .clk(clk),
      .out(par_done_reg692_out),
      .done(par_done_reg692_done)
  );
  
  std_reg #(1) par_done_reg693 (
      .in(par_done_reg693_in),
      .write_en(par_done_reg693_write_en),
      .clk(clk),
      .out(par_done_reg693_out),
      .done(par_done_reg693_done)
  );
  
  std_reg #(1) par_done_reg694 (
      .in(par_done_reg694_in),
      .write_en(par_done_reg694_write_en),
      .clk(clk),
      .out(par_done_reg694_out),
      .done(par_done_reg694_done)
  );
  
  std_reg #(1) par_done_reg695 (
      .in(par_done_reg695_in),
      .write_en(par_done_reg695_write_en),
      .clk(clk),
      .out(par_done_reg695_out),
      .done(par_done_reg695_done)
  );
  
  std_reg #(1) par_done_reg696 (
      .in(par_done_reg696_in),
      .write_en(par_done_reg696_write_en),
      .clk(clk),
      .out(par_done_reg696_out),
      .done(par_done_reg696_done)
  );
  
  std_reg #(1) par_done_reg697 (
      .in(par_done_reg697_in),
      .write_en(par_done_reg697_write_en),
      .clk(clk),
      .out(par_done_reg697_out),
      .done(par_done_reg697_done)
  );
  
  std_reg #(1) par_done_reg698 (
      .in(par_done_reg698_in),
      .write_en(par_done_reg698_write_en),
      .clk(clk),
      .out(par_done_reg698_out),
      .done(par_done_reg698_done)
  );
  
  std_reg #(1) par_done_reg699 (
      .in(par_done_reg699_in),
      .write_en(par_done_reg699_write_en),
      .clk(clk),
      .out(par_done_reg699_out),
      .done(par_done_reg699_done)
  );
  
  std_reg #(1) par_done_reg700 (
      .in(par_done_reg700_in),
      .write_en(par_done_reg700_write_en),
      .clk(clk),
      .out(par_done_reg700_out),
      .done(par_done_reg700_done)
  );
  
  std_reg #(1) par_done_reg701 (
      .in(par_done_reg701_in),
      .write_en(par_done_reg701_write_en),
      .clk(clk),
      .out(par_done_reg701_out),
      .done(par_done_reg701_done)
  );
  
  std_reg #(1) par_done_reg702 (
      .in(par_done_reg702_in),
      .write_en(par_done_reg702_write_en),
      .clk(clk),
      .out(par_done_reg702_out),
      .done(par_done_reg702_done)
  );
  
  std_reg #(1) par_done_reg703 (
      .in(par_done_reg703_in),
      .write_en(par_done_reg703_write_en),
      .clk(clk),
      .out(par_done_reg703_out),
      .done(par_done_reg703_done)
  );
  
  std_reg #(1) par_done_reg704 (
      .in(par_done_reg704_in),
      .write_en(par_done_reg704_write_en),
      .clk(clk),
      .out(par_done_reg704_out),
      .done(par_done_reg704_done)
  );
  
  std_reg #(1) par_done_reg705 (
      .in(par_done_reg705_in),
      .write_en(par_done_reg705_write_en),
      .clk(clk),
      .out(par_done_reg705_out),
      .done(par_done_reg705_done)
  );
  
  std_reg #(1) par_done_reg706 (
      .in(par_done_reg706_in),
      .write_en(par_done_reg706_write_en),
      .clk(clk),
      .out(par_done_reg706_out),
      .done(par_done_reg706_done)
  );
  
  std_reg #(1) par_done_reg707 (
      .in(par_done_reg707_in),
      .write_en(par_done_reg707_write_en),
      .clk(clk),
      .out(par_done_reg707_out),
      .done(par_done_reg707_done)
  );
  
  std_reg #(1) par_done_reg708 (
      .in(par_done_reg708_in),
      .write_en(par_done_reg708_write_en),
      .clk(clk),
      .out(par_done_reg708_out),
      .done(par_done_reg708_done)
  );
  
  std_reg #(1) par_done_reg709 (
      .in(par_done_reg709_in),
      .write_en(par_done_reg709_write_en),
      .clk(clk),
      .out(par_done_reg709_out),
      .done(par_done_reg709_done)
  );
  
  std_reg #(1) par_done_reg710 (
      .in(par_done_reg710_in),
      .write_en(par_done_reg710_write_en),
      .clk(clk),
      .out(par_done_reg710_out),
      .done(par_done_reg710_done)
  );
  
  std_reg #(1) par_done_reg711 (
      .in(par_done_reg711_in),
      .write_en(par_done_reg711_write_en),
      .clk(clk),
      .out(par_done_reg711_out),
      .done(par_done_reg711_done)
  );
  
  std_reg #(1) par_done_reg712 (
      .in(par_done_reg712_in),
      .write_en(par_done_reg712_write_en),
      .clk(clk),
      .out(par_done_reg712_out),
      .done(par_done_reg712_done)
  );
  
  std_reg #(1) par_done_reg713 (
      .in(par_done_reg713_in),
      .write_en(par_done_reg713_write_en),
      .clk(clk),
      .out(par_done_reg713_out),
      .done(par_done_reg713_done)
  );
  
  std_reg #(1) par_done_reg714 (
      .in(par_done_reg714_in),
      .write_en(par_done_reg714_write_en),
      .clk(clk),
      .out(par_done_reg714_out),
      .done(par_done_reg714_done)
  );
  
  std_reg #(1) par_done_reg715 (
      .in(par_done_reg715_in),
      .write_en(par_done_reg715_write_en),
      .clk(clk),
      .out(par_done_reg715_out),
      .done(par_done_reg715_done)
  );
  
  std_reg #(1) par_done_reg716 (
      .in(par_done_reg716_in),
      .write_en(par_done_reg716_write_en),
      .clk(clk),
      .out(par_done_reg716_out),
      .done(par_done_reg716_done)
  );
  
  std_reg #(1) par_done_reg717 (
      .in(par_done_reg717_in),
      .write_en(par_done_reg717_write_en),
      .clk(clk),
      .out(par_done_reg717_out),
      .done(par_done_reg717_done)
  );
  
  std_reg #(1) par_done_reg718 (
      .in(par_done_reg718_in),
      .write_en(par_done_reg718_write_en),
      .clk(clk),
      .out(par_done_reg718_out),
      .done(par_done_reg718_done)
  );
  
  std_reg #(1) par_done_reg719 (
      .in(par_done_reg719_in),
      .write_en(par_done_reg719_write_en),
      .clk(clk),
      .out(par_done_reg719_out),
      .done(par_done_reg719_done)
  );
  
  std_reg #(1) par_done_reg720 (
      .in(par_done_reg720_in),
      .write_en(par_done_reg720_write_en),
      .clk(clk),
      .out(par_done_reg720_out),
      .done(par_done_reg720_done)
  );
  
  std_reg #(1) par_done_reg721 (
      .in(par_done_reg721_in),
      .write_en(par_done_reg721_write_en),
      .clk(clk),
      .out(par_done_reg721_out),
      .done(par_done_reg721_done)
  );
  
  std_reg #(1) par_done_reg722 (
      .in(par_done_reg722_in),
      .write_en(par_done_reg722_write_en),
      .clk(clk),
      .out(par_done_reg722_out),
      .done(par_done_reg722_done)
  );
  
  std_reg #(1) par_done_reg723 (
      .in(par_done_reg723_in),
      .write_en(par_done_reg723_write_en),
      .clk(clk),
      .out(par_done_reg723_out),
      .done(par_done_reg723_done)
  );
  
  std_reg #(1) par_done_reg724 (
      .in(par_done_reg724_in),
      .write_en(par_done_reg724_write_en),
      .clk(clk),
      .out(par_done_reg724_out),
      .done(par_done_reg724_done)
  );
  
  std_reg #(1) par_done_reg725 (
      .in(par_done_reg725_in),
      .write_en(par_done_reg725_write_en),
      .clk(clk),
      .out(par_done_reg725_out),
      .done(par_done_reg725_done)
  );
  
  std_reg #(1) par_done_reg726 (
      .in(par_done_reg726_in),
      .write_en(par_done_reg726_write_en),
      .clk(clk),
      .out(par_done_reg726_out),
      .done(par_done_reg726_done)
  );
  
  std_reg #(1) par_done_reg727 (
      .in(par_done_reg727_in),
      .write_en(par_done_reg727_write_en),
      .clk(clk),
      .out(par_done_reg727_out),
      .done(par_done_reg727_done)
  );
  
  std_reg #(1) par_done_reg728 (
      .in(par_done_reg728_in),
      .write_en(par_done_reg728_write_en),
      .clk(clk),
      .out(par_done_reg728_out),
      .done(par_done_reg728_done)
  );
  
  std_reg #(1) par_done_reg729 (
      .in(par_done_reg729_in),
      .write_en(par_done_reg729_write_en),
      .clk(clk),
      .out(par_done_reg729_out),
      .done(par_done_reg729_done)
  );
  
  std_reg #(1) par_done_reg730 (
      .in(par_done_reg730_in),
      .write_en(par_done_reg730_write_en),
      .clk(clk),
      .out(par_done_reg730_out),
      .done(par_done_reg730_done)
  );
  
  std_reg #(1) par_done_reg731 (
      .in(par_done_reg731_in),
      .write_en(par_done_reg731_write_en),
      .clk(clk),
      .out(par_done_reg731_out),
      .done(par_done_reg731_done)
  );
  
  std_reg #(1) par_done_reg732 (
      .in(par_done_reg732_in),
      .write_en(par_done_reg732_write_en),
      .clk(clk),
      .out(par_done_reg732_out),
      .done(par_done_reg732_done)
  );
  
  std_reg #(1) par_done_reg733 (
      .in(par_done_reg733_in),
      .write_en(par_done_reg733_write_en),
      .clk(clk),
      .out(par_done_reg733_out),
      .done(par_done_reg733_done)
  );
  
  std_reg #(1) par_done_reg734 (
      .in(par_done_reg734_in),
      .write_en(par_done_reg734_write_en),
      .clk(clk),
      .out(par_done_reg734_out),
      .done(par_done_reg734_done)
  );
  
  std_reg #(1) par_done_reg735 (
      .in(par_done_reg735_in),
      .write_en(par_done_reg735_write_en),
      .clk(clk),
      .out(par_done_reg735_out),
      .done(par_done_reg735_done)
  );
  
  std_reg #(1) par_done_reg736 (
      .in(par_done_reg736_in),
      .write_en(par_done_reg736_write_en),
      .clk(clk),
      .out(par_done_reg736_out),
      .done(par_done_reg736_done)
  );
  
  std_reg #(1) par_done_reg737 (
      .in(par_done_reg737_in),
      .write_en(par_done_reg737_write_en),
      .clk(clk),
      .out(par_done_reg737_out),
      .done(par_done_reg737_done)
  );
  
  std_reg #(1) par_done_reg738 (
      .in(par_done_reg738_in),
      .write_en(par_done_reg738_write_en),
      .clk(clk),
      .out(par_done_reg738_out),
      .done(par_done_reg738_done)
  );
  
  std_reg #(1) par_done_reg739 (
      .in(par_done_reg739_in),
      .write_en(par_done_reg739_write_en),
      .clk(clk),
      .out(par_done_reg739_out),
      .done(par_done_reg739_done)
  );
  
  std_reg #(1) par_done_reg740 (
      .in(par_done_reg740_in),
      .write_en(par_done_reg740_write_en),
      .clk(clk),
      .out(par_done_reg740_out),
      .done(par_done_reg740_done)
  );
  
  std_reg #(1) par_done_reg741 (
      .in(par_done_reg741_in),
      .write_en(par_done_reg741_write_en),
      .clk(clk),
      .out(par_done_reg741_out),
      .done(par_done_reg741_done)
  );
  
  std_reg #(1) par_done_reg742 (
      .in(par_done_reg742_in),
      .write_en(par_done_reg742_write_en),
      .clk(clk),
      .out(par_done_reg742_out),
      .done(par_done_reg742_done)
  );
  
  std_reg #(1) par_done_reg743 (
      .in(par_done_reg743_in),
      .write_en(par_done_reg743_write_en),
      .clk(clk),
      .out(par_done_reg743_out),
      .done(par_done_reg743_done)
  );
  
  std_reg #(1) par_done_reg744 (
      .in(par_done_reg744_in),
      .write_en(par_done_reg744_write_en),
      .clk(clk),
      .out(par_done_reg744_out),
      .done(par_done_reg744_done)
  );
  
  std_reg #(1) par_done_reg745 (
      .in(par_done_reg745_in),
      .write_en(par_done_reg745_write_en),
      .clk(clk),
      .out(par_done_reg745_out),
      .done(par_done_reg745_done)
  );
  
  std_reg #(1) par_done_reg746 (
      .in(par_done_reg746_in),
      .write_en(par_done_reg746_write_en),
      .clk(clk),
      .out(par_done_reg746_out),
      .done(par_done_reg746_done)
  );
  
  std_reg #(1) par_done_reg747 (
      .in(par_done_reg747_in),
      .write_en(par_done_reg747_write_en),
      .clk(clk),
      .out(par_done_reg747_out),
      .done(par_done_reg747_done)
  );
  
  std_reg #(1) par_reset22 (
      .in(par_reset22_in),
      .write_en(par_reset22_write_en),
      .clk(clk),
      .out(par_reset22_out),
      .done(par_reset22_done)
  );
  
  std_reg #(1) par_done_reg748 (
      .in(par_done_reg748_in),
      .write_en(par_done_reg748_write_en),
      .clk(clk),
      .out(par_done_reg748_out),
      .done(par_done_reg748_done)
  );
  
  std_reg #(1) par_done_reg749 (
      .in(par_done_reg749_in),
      .write_en(par_done_reg749_write_en),
      .clk(clk),
      .out(par_done_reg749_out),
      .done(par_done_reg749_done)
  );
  
  std_reg #(1) par_done_reg750 (
      .in(par_done_reg750_in),
      .write_en(par_done_reg750_write_en),
      .clk(clk),
      .out(par_done_reg750_out),
      .done(par_done_reg750_done)
  );
  
  std_reg #(1) par_done_reg751 (
      .in(par_done_reg751_in),
      .write_en(par_done_reg751_write_en),
      .clk(clk),
      .out(par_done_reg751_out),
      .done(par_done_reg751_done)
  );
  
  std_reg #(1) par_done_reg752 (
      .in(par_done_reg752_in),
      .write_en(par_done_reg752_write_en),
      .clk(clk),
      .out(par_done_reg752_out),
      .done(par_done_reg752_done)
  );
  
  std_reg #(1) par_done_reg753 (
      .in(par_done_reg753_in),
      .write_en(par_done_reg753_write_en),
      .clk(clk),
      .out(par_done_reg753_out),
      .done(par_done_reg753_done)
  );
  
  std_reg #(1) par_done_reg754 (
      .in(par_done_reg754_in),
      .write_en(par_done_reg754_write_en),
      .clk(clk),
      .out(par_done_reg754_out),
      .done(par_done_reg754_done)
  );
  
  std_reg #(1) par_done_reg755 (
      .in(par_done_reg755_in),
      .write_en(par_done_reg755_write_en),
      .clk(clk),
      .out(par_done_reg755_out),
      .done(par_done_reg755_done)
  );
  
  std_reg #(1) par_done_reg756 (
      .in(par_done_reg756_in),
      .write_en(par_done_reg756_write_en),
      .clk(clk),
      .out(par_done_reg756_out),
      .done(par_done_reg756_done)
  );
  
  std_reg #(1) par_done_reg757 (
      .in(par_done_reg757_in),
      .write_en(par_done_reg757_write_en),
      .clk(clk),
      .out(par_done_reg757_out),
      .done(par_done_reg757_done)
  );
  
  std_reg #(1) par_done_reg758 (
      .in(par_done_reg758_in),
      .write_en(par_done_reg758_write_en),
      .clk(clk),
      .out(par_done_reg758_out),
      .done(par_done_reg758_done)
  );
  
  std_reg #(1) par_done_reg759 (
      .in(par_done_reg759_in),
      .write_en(par_done_reg759_write_en),
      .clk(clk),
      .out(par_done_reg759_out),
      .done(par_done_reg759_done)
  );
  
  std_reg #(1) par_done_reg760 (
      .in(par_done_reg760_in),
      .write_en(par_done_reg760_write_en),
      .clk(clk),
      .out(par_done_reg760_out),
      .done(par_done_reg760_done)
  );
  
  std_reg #(1) par_done_reg761 (
      .in(par_done_reg761_in),
      .write_en(par_done_reg761_write_en),
      .clk(clk),
      .out(par_done_reg761_out),
      .done(par_done_reg761_done)
  );
  
  std_reg #(1) par_done_reg762 (
      .in(par_done_reg762_in),
      .write_en(par_done_reg762_write_en),
      .clk(clk),
      .out(par_done_reg762_out),
      .done(par_done_reg762_done)
  );
  
  std_reg #(1) par_done_reg763 (
      .in(par_done_reg763_in),
      .write_en(par_done_reg763_write_en),
      .clk(clk),
      .out(par_done_reg763_out),
      .done(par_done_reg763_done)
  );
  
  std_reg #(1) par_done_reg764 (
      .in(par_done_reg764_in),
      .write_en(par_done_reg764_write_en),
      .clk(clk),
      .out(par_done_reg764_out),
      .done(par_done_reg764_done)
  );
  
  std_reg #(1) par_done_reg765 (
      .in(par_done_reg765_in),
      .write_en(par_done_reg765_write_en),
      .clk(clk),
      .out(par_done_reg765_out),
      .done(par_done_reg765_done)
  );
  
  std_reg #(1) par_done_reg766 (
      .in(par_done_reg766_in),
      .write_en(par_done_reg766_write_en),
      .clk(clk),
      .out(par_done_reg766_out),
      .done(par_done_reg766_done)
  );
  
  std_reg #(1) par_done_reg767 (
      .in(par_done_reg767_in),
      .write_en(par_done_reg767_write_en),
      .clk(clk),
      .out(par_done_reg767_out),
      .done(par_done_reg767_done)
  );
  
  std_reg #(1) par_done_reg768 (
      .in(par_done_reg768_in),
      .write_en(par_done_reg768_write_en),
      .clk(clk),
      .out(par_done_reg768_out),
      .done(par_done_reg768_done)
  );
  
  std_reg #(1) par_done_reg769 (
      .in(par_done_reg769_in),
      .write_en(par_done_reg769_write_en),
      .clk(clk),
      .out(par_done_reg769_out),
      .done(par_done_reg769_done)
  );
  
  std_reg #(1) par_done_reg770 (
      .in(par_done_reg770_in),
      .write_en(par_done_reg770_write_en),
      .clk(clk),
      .out(par_done_reg770_out),
      .done(par_done_reg770_done)
  );
  
  std_reg #(1) par_done_reg771 (
      .in(par_done_reg771_in),
      .write_en(par_done_reg771_write_en),
      .clk(clk),
      .out(par_done_reg771_out),
      .done(par_done_reg771_done)
  );
  
  std_reg #(1) par_done_reg772 (
      .in(par_done_reg772_in),
      .write_en(par_done_reg772_write_en),
      .clk(clk),
      .out(par_done_reg772_out),
      .done(par_done_reg772_done)
  );
  
  std_reg #(1) par_done_reg773 (
      .in(par_done_reg773_in),
      .write_en(par_done_reg773_write_en),
      .clk(clk),
      .out(par_done_reg773_out),
      .done(par_done_reg773_done)
  );
  
  std_reg #(1) par_done_reg774 (
      .in(par_done_reg774_in),
      .write_en(par_done_reg774_write_en),
      .clk(clk),
      .out(par_done_reg774_out),
      .done(par_done_reg774_done)
  );
  
  std_reg #(1) par_done_reg775 (
      .in(par_done_reg775_in),
      .write_en(par_done_reg775_write_en),
      .clk(clk),
      .out(par_done_reg775_out),
      .done(par_done_reg775_done)
  );
  
  std_reg #(1) par_done_reg776 (
      .in(par_done_reg776_in),
      .write_en(par_done_reg776_write_en),
      .clk(clk),
      .out(par_done_reg776_out),
      .done(par_done_reg776_done)
  );
  
  std_reg #(1) par_done_reg777 (
      .in(par_done_reg777_in),
      .write_en(par_done_reg777_write_en),
      .clk(clk),
      .out(par_done_reg777_out),
      .done(par_done_reg777_done)
  );
  
  std_reg #(1) par_done_reg778 (
      .in(par_done_reg778_in),
      .write_en(par_done_reg778_write_en),
      .clk(clk),
      .out(par_done_reg778_out),
      .done(par_done_reg778_done)
  );
  
  std_reg #(1) par_done_reg779 (
      .in(par_done_reg779_in),
      .write_en(par_done_reg779_write_en),
      .clk(clk),
      .out(par_done_reg779_out),
      .done(par_done_reg779_done)
  );
  
  std_reg #(1) par_done_reg780 (
      .in(par_done_reg780_in),
      .write_en(par_done_reg780_write_en),
      .clk(clk),
      .out(par_done_reg780_out),
      .done(par_done_reg780_done)
  );
  
  std_reg #(1) par_done_reg781 (
      .in(par_done_reg781_in),
      .write_en(par_done_reg781_write_en),
      .clk(clk),
      .out(par_done_reg781_out),
      .done(par_done_reg781_done)
  );
  
  std_reg #(1) par_done_reg782 (
      .in(par_done_reg782_in),
      .write_en(par_done_reg782_write_en),
      .clk(clk),
      .out(par_done_reg782_out),
      .done(par_done_reg782_done)
  );
  
  std_reg #(1) par_done_reg783 (
      .in(par_done_reg783_in),
      .write_en(par_done_reg783_write_en),
      .clk(clk),
      .out(par_done_reg783_out),
      .done(par_done_reg783_done)
  );
  
  std_reg #(1) par_done_reg784 (
      .in(par_done_reg784_in),
      .write_en(par_done_reg784_write_en),
      .clk(clk),
      .out(par_done_reg784_out),
      .done(par_done_reg784_done)
  );
  
  std_reg #(1) par_done_reg785 (
      .in(par_done_reg785_in),
      .write_en(par_done_reg785_write_en),
      .clk(clk),
      .out(par_done_reg785_out),
      .done(par_done_reg785_done)
  );
  
  std_reg #(1) par_done_reg786 (
      .in(par_done_reg786_in),
      .write_en(par_done_reg786_write_en),
      .clk(clk),
      .out(par_done_reg786_out),
      .done(par_done_reg786_done)
  );
  
  std_reg #(1) par_done_reg787 (
      .in(par_done_reg787_in),
      .write_en(par_done_reg787_write_en),
      .clk(clk),
      .out(par_done_reg787_out),
      .done(par_done_reg787_done)
  );
  
  std_reg #(1) par_done_reg788 (
      .in(par_done_reg788_in),
      .write_en(par_done_reg788_write_en),
      .clk(clk),
      .out(par_done_reg788_out),
      .done(par_done_reg788_done)
  );
  
  std_reg #(1) par_done_reg789 (
      .in(par_done_reg789_in),
      .write_en(par_done_reg789_write_en),
      .clk(clk),
      .out(par_done_reg789_out),
      .done(par_done_reg789_done)
  );
  
  std_reg #(1) par_done_reg790 (
      .in(par_done_reg790_in),
      .write_en(par_done_reg790_write_en),
      .clk(clk),
      .out(par_done_reg790_out),
      .done(par_done_reg790_done)
  );
  
  std_reg #(1) par_done_reg791 (
      .in(par_done_reg791_in),
      .write_en(par_done_reg791_write_en),
      .clk(clk),
      .out(par_done_reg791_out),
      .done(par_done_reg791_done)
  );
  
  std_reg #(1) par_done_reg792 (
      .in(par_done_reg792_in),
      .write_en(par_done_reg792_write_en),
      .clk(clk),
      .out(par_done_reg792_out),
      .done(par_done_reg792_done)
  );
  
  std_reg #(1) par_done_reg793 (
      .in(par_done_reg793_in),
      .write_en(par_done_reg793_write_en),
      .clk(clk),
      .out(par_done_reg793_out),
      .done(par_done_reg793_done)
  );
  
  std_reg #(1) par_done_reg794 (
      .in(par_done_reg794_in),
      .write_en(par_done_reg794_write_en),
      .clk(clk),
      .out(par_done_reg794_out),
      .done(par_done_reg794_done)
  );
  
  std_reg #(1) par_done_reg795 (
      .in(par_done_reg795_in),
      .write_en(par_done_reg795_write_en),
      .clk(clk),
      .out(par_done_reg795_out),
      .done(par_done_reg795_done)
  );
  
  std_reg #(1) par_done_reg796 (
      .in(par_done_reg796_in),
      .write_en(par_done_reg796_write_en),
      .clk(clk),
      .out(par_done_reg796_out),
      .done(par_done_reg796_done)
  );
  
  std_reg #(1) par_done_reg797 (
      .in(par_done_reg797_in),
      .write_en(par_done_reg797_write_en),
      .clk(clk),
      .out(par_done_reg797_out),
      .done(par_done_reg797_done)
  );
  
  std_reg #(1) par_done_reg798 (
      .in(par_done_reg798_in),
      .write_en(par_done_reg798_write_en),
      .clk(clk),
      .out(par_done_reg798_out),
      .done(par_done_reg798_done)
  );
  
  std_reg #(1) par_done_reg799 (
      .in(par_done_reg799_in),
      .write_en(par_done_reg799_write_en),
      .clk(clk),
      .out(par_done_reg799_out),
      .done(par_done_reg799_done)
  );
  
  std_reg #(1) par_done_reg800 (
      .in(par_done_reg800_in),
      .write_en(par_done_reg800_write_en),
      .clk(clk),
      .out(par_done_reg800_out),
      .done(par_done_reg800_done)
  );
  
  std_reg #(1) par_done_reg801 (
      .in(par_done_reg801_in),
      .write_en(par_done_reg801_write_en),
      .clk(clk),
      .out(par_done_reg801_out),
      .done(par_done_reg801_done)
  );
  
  std_reg #(1) par_done_reg802 (
      .in(par_done_reg802_in),
      .write_en(par_done_reg802_write_en),
      .clk(clk),
      .out(par_done_reg802_out),
      .done(par_done_reg802_done)
  );
  
  std_reg #(1) par_done_reg803 (
      .in(par_done_reg803_in),
      .write_en(par_done_reg803_write_en),
      .clk(clk),
      .out(par_done_reg803_out),
      .done(par_done_reg803_done)
  );
  
  std_reg #(1) par_done_reg804 (
      .in(par_done_reg804_in),
      .write_en(par_done_reg804_write_en),
      .clk(clk),
      .out(par_done_reg804_out),
      .done(par_done_reg804_done)
  );
  
  std_reg #(1) par_done_reg805 (
      .in(par_done_reg805_in),
      .write_en(par_done_reg805_write_en),
      .clk(clk),
      .out(par_done_reg805_out),
      .done(par_done_reg805_done)
  );
  
  std_reg #(1) par_done_reg806 (
      .in(par_done_reg806_in),
      .write_en(par_done_reg806_write_en),
      .clk(clk),
      .out(par_done_reg806_out),
      .done(par_done_reg806_done)
  );
  
  std_reg #(1) par_done_reg807 (
      .in(par_done_reg807_in),
      .write_en(par_done_reg807_write_en),
      .clk(clk),
      .out(par_done_reg807_out),
      .done(par_done_reg807_done)
  );
  
  std_reg #(1) par_done_reg808 (
      .in(par_done_reg808_in),
      .write_en(par_done_reg808_write_en),
      .clk(clk),
      .out(par_done_reg808_out),
      .done(par_done_reg808_done)
  );
  
  std_reg #(1) par_done_reg809 (
      .in(par_done_reg809_in),
      .write_en(par_done_reg809_write_en),
      .clk(clk),
      .out(par_done_reg809_out),
      .done(par_done_reg809_done)
  );
  
  std_reg #(1) par_done_reg810 (
      .in(par_done_reg810_in),
      .write_en(par_done_reg810_write_en),
      .clk(clk),
      .out(par_done_reg810_out),
      .done(par_done_reg810_done)
  );
  
  std_reg #(1) par_done_reg811 (
      .in(par_done_reg811_in),
      .write_en(par_done_reg811_write_en),
      .clk(clk),
      .out(par_done_reg811_out),
      .done(par_done_reg811_done)
  );
  
  std_reg #(1) par_done_reg812 (
      .in(par_done_reg812_in),
      .write_en(par_done_reg812_write_en),
      .clk(clk),
      .out(par_done_reg812_out),
      .done(par_done_reg812_done)
  );
  
  std_reg #(1) par_done_reg813 (
      .in(par_done_reg813_in),
      .write_en(par_done_reg813_write_en),
      .clk(clk),
      .out(par_done_reg813_out),
      .done(par_done_reg813_done)
  );
  
  std_reg #(1) par_done_reg814 (
      .in(par_done_reg814_in),
      .write_en(par_done_reg814_write_en),
      .clk(clk),
      .out(par_done_reg814_out),
      .done(par_done_reg814_done)
  );
  
  std_reg #(1) par_done_reg815 (
      .in(par_done_reg815_in),
      .write_en(par_done_reg815_write_en),
      .clk(clk),
      .out(par_done_reg815_out),
      .done(par_done_reg815_done)
  );
  
  std_reg #(1) par_done_reg816 (
      .in(par_done_reg816_in),
      .write_en(par_done_reg816_write_en),
      .clk(clk),
      .out(par_done_reg816_out),
      .done(par_done_reg816_done)
  );
  
  std_reg #(1) par_done_reg817 (
      .in(par_done_reg817_in),
      .write_en(par_done_reg817_write_en),
      .clk(clk),
      .out(par_done_reg817_out),
      .done(par_done_reg817_done)
  );
  
  std_reg #(1) par_done_reg818 (
      .in(par_done_reg818_in),
      .write_en(par_done_reg818_write_en),
      .clk(clk),
      .out(par_done_reg818_out),
      .done(par_done_reg818_done)
  );
  
  std_reg #(1) par_done_reg819 (
      .in(par_done_reg819_in),
      .write_en(par_done_reg819_write_en),
      .clk(clk),
      .out(par_done_reg819_out),
      .done(par_done_reg819_done)
  );
  
  std_reg #(1) par_done_reg820 (
      .in(par_done_reg820_in),
      .write_en(par_done_reg820_write_en),
      .clk(clk),
      .out(par_done_reg820_out),
      .done(par_done_reg820_done)
  );
  
  std_reg #(1) par_done_reg821 (
      .in(par_done_reg821_in),
      .write_en(par_done_reg821_write_en),
      .clk(clk),
      .out(par_done_reg821_out),
      .done(par_done_reg821_done)
  );
  
  std_reg #(1) par_done_reg822 (
      .in(par_done_reg822_in),
      .write_en(par_done_reg822_write_en),
      .clk(clk),
      .out(par_done_reg822_out),
      .done(par_done_reg822_done)
  );
  
  std_reg #(1) par_done_reg823 (
      .in(par_done_reg823_in),
      .write_en(par_done_reg823_write_en),
      .clk(clk),
      .out(par_done_reg823_out),
      .done(par_done_reg823_done)
  );
  
  std_reg #(1) par_done_reg824 (
      .in(par_done_reg824_in),
      .write_en(par_done_reg824_write_en),
      .clk(clk),
      .out(par_done_reg824_out),
      .done(par_done_reg824_done)
  );
  
  std_reg #(1) par_done_reg825 (
      .in(par_done_reg825_in),
      .write_en(par_done_reg825_write_en),
      .clk(clk),
      .out(par_done_reg825_out),
      .done(par_done_reg825_done)
  );
  
  std_reg #(1) par_done_reg826 (
      .in(par_done_reg826_in),
      .write_en(par_done_reg826_write_en),
      .clk(clk),
      .out(par_done_reg826_out),
      .done(par_done_reg826_done)
  );
  
  std_reg #(1) par_done_reg827 (
      .in(par_done_reg827_in),
      .write_en(par_done_reg827_write_en),
      .clk(clk),
      .out(par_done_reg827_out),
      .done(par_done_reg827_done)
  );
  
  std_reg #(1) par_done_reg828 (
      .in(par_done_reg828_in),
      .write_en(par_done_reg828_write_en),
      .clk(clk),
      .out(par_done_reg828_out),
      .done(par_done_reg828_done)
  );
  
  std_reg #(1) par_done_reg829 (
      .in(par_done_reg829_in),
      .write_en(par_done_reg829_write_en),
      .clk(clk),
      .out(par_done_reg829_out),
      .done(par_done_reg829_done)
  );
  
  std_reg #(1) par_done_reg830 (
      .in(par_done_reg830_in),
      .write_en(par_done_reg830_write_en),
      .clk(clk),
      .out(par_done_reg830_out),
      .done(par_done_reg830_done)
  );
  
  std_reg #(1) par_done_reg831 (
      .in(par_done_reg831_in),
      .write_en(par_done_reg831_write_en),
      .clk(clk),
      .out(par_done_reg831_out),
      .done(par_done_reg831_done)
  );
  
  std_reg #(1) par_done_reg832 (
      .in(par_done_reg832_in),
      .write_en(par_done_reg832_write_en),
      .clk(clk),
      .out(par_done_reg832_out),
      .done(par_done_reg832_done)
  );
  
  std_reg #(1) par_done_reg833 (
      .in(par_done_reg833_in),
      .write_en(par_done_reg833_write_en),
      .clk(clk),
      .out(par_done_reg833_out),
      .done(par_done_reg833_done)
  );
  
  std_reg #(1) par_done_reg834 (
      .in(par_done_reg834_in),
      .write_en(par_done_reg834_write_en),
      .clk(clk),
      .out(par_done_reg834_out),
      .done(par_done_reg834_done)
  );
  
  std_reg #(1) par_done_reg835 (
      .in(par_done_reg835_in),
      .write_en(par_done_reg835_write_en),
      .clk(clk),
      .out(par_done_reg835_out),
      .done(par_done_reg835_done)
  );
  
  std_reg #(1) par_done_reg836 (
      .in(par_done_reg836_in),
      .write_en(par_done_reg836_write_en),
      .clk(clk),
      .out(par_done_reg836_out),
      .done(par_done_reg836_done)
  );
  
  std_reg #(1) par_done_reg837 (
      .in(par_done_reg837_in),
      .write_en(par_done_reg837_write_en),
      .clk(clk),
      .out(par_done_reg837_out),
      .done(par_done_reg837_done)
  );
  
  std_reg #(1) par_done_reg838 (
      .in(par_done_reg838_in),
      .write_en(par_done_reg838_write_en),
      .clk(clk),
      .out(par_done_reg838_out),
      .done(par_done_reg838_done)
  );
  
  std_reg #(1) par_done_reg839 (
      .in(par_done_reg839_in),
      .write_en(par_done_reg839_write_en),
      .clk(clk),
      .out(par_done_reg839_out),
      .done(par_done_reg839_done)
  );
  
  std_reg #(1) par_done_reg840 (
      .in(par_done_reg840_in),
      .write_en(par_done_reg840_write_en),
      .clk(clk),
      .out(par_done_reg840_out),
      .done(par_done_reg840_done)
  );
  
  std_reg #(1) par_done_reg841 (
      .in(par_done_reg841_in),
      .write_en(par_done_reg841_write_en),
      .clk(clk),
      .out(par_done_reg841_out),
      .done(par_done_reg841_done)
  );
  
  std_reg #(1) par_done_reg842 (
      .in(par_done_reg842_in),
      .write_en(par_done_reg842_write_en),
      .clk(clk),
      .out(par_done_reg842_out),
      .done(par_done_reg842_done)
  );
  
  std_reg #(1) par_done_reg843 (
      .in(par_done_reg843_in),
      .write_en(par_done_reg843_write_en),
      .clk(clk),
      .out(par_done_reg843_out),
      .done(par_done_reg843_done)
  );
  
  std_reg #(1) par_reset23 (
      .in(par_reset23_in),
      .write_en(par_reset23_write_en),
      .clk(clk),
      .out(par_reset23_out),
      .done(par_reset23_done)
  );
  
  std_reg #(1) par_done_reg844 (
      .in(par_done_reg844_in),
      .write_en(par_done_reg844_write_en),
      .clk(clk),
      .out(par_done_reg844_out),
      .done(par_done_reg844_done)
  );
  
  std_reg #(1) par_done_reg845 (
      .in(par_done_reg845_in),
      .write_en(par_done_reg845_write_en),
      .clk(clk),
      .out(par_done_reg845_out),
      .done(par_done_reg845_done)
  );
  
  std_reg #(1) par_done_reg846 (
      .in(par_done_reg846_in),
      .write_en(par_done_reg846_write_en),
      .clk(clk),
      .out(par_done_reg846_out),
      .done(par_done_reg846_done)
  );
  
  std_reg #(1) par_done_reg847 (
      .in(par_done_reg847_in),
      .write_en(par_done_reg847_write_en),
      .clk(clk),
      .out(par_done_reg847_out),
      .done(par_done_reg847_done)
  );
  
  std_reg #(1) par_done_reg848 (
      .in(par_done_reg848_in),
      .write_en(par_done_reg848_write_en),
      .clk(clk),
      .out(par_done_reg848_out),
      .done(par_done_reg848_done)
  );
  
  std_reg #(1) par_done_reg849 (
      .in(par_done_reg849_in),
      .write_en(par_done_reg849_write_en),
      .clk(clk),
      .out(par_done_reg849_out),
      .done(par_done_reg849_done)
  );
  
  std_reg #(1) par_done_reg850 (
      .in(par_done_reg850_in),
      .write_en(par_done_reg850_write_en),
      .clk(clk),
      .out(par_done_reg850_out),
      .done(par_done_reg850_done)
  );
  
  std_reg #(1) par_done_reg851 (
      .in(par_done_reg851_in),
      .write_en(par_done_reg851_write_en),
      .clk(clk),
      .out(par_done_reg851_out),
      .done(par_done_reg851_done)
  );
  
  std_reg #(1) par_done_reg852 (
      .in(par_done_reg852_in),
      .write_en(par_done_reg852_write_en),
      .clk(clk),
      .out(par_done_reg852_out),
      .done(par_done_reg852_done)
  );
  
  std_reg #(1) par_done_reg853 (
      .in(par_done_reg853_in),
      .write_en(par_done_reg853_write_en),
      .clk(clk),
      .out(par_done_reg853_out),
      .done(par_done_reg853_done)
  );
  
  std_reg #(1) par_done_reg854 (
      .in(par_done_reg854_in),
      .write_en(par_done_reg854_write_en),
      .clk(clk),
      .out(par_done_reg854_out),
      .done(par_done_reg854_done)
  );
  
  std_reg #(1) par_done_reg855 (
      .in(par_done_reg855_in),
      .write_en(par_done_reg855_write_en),
      .clk(clk),
      .out(par_done_reg855_out),
      .done(par_done_reg855_done)
  );
  
  std_reg #(1) par_done_reg856 (
      .in(par_done_reg856_in),
      .write_en(par_done_reg856_write_en),
      .clk(clk),
      .out(par_done_reg856_out),
      .done(par_done_reg856_done)
  );
  
  std_reg #(1) par_done_reg857 (
      .in(par_done_reg857_in),
      .write_en(par_done_reg857_write_en),
      .clk(clk),
      .out(par_done_reg857_out),
      .done(par_done_reg857_done)
  );
  
  std_reg #(1) par_done_reg858 (
      .in(par_done_reg858_in),
      .write_en(par_done_reg858_write_en),
      .clk(clk),
      .out(par_done_reg858_out),
      .done(par_done_reg858_done)
  );
  
  std_reg #(1) par_done_reg859 (
      .in(par_done_reg859_in),
      .write_en(par_done_reg859_write_en),
      .clk(clk),
      .out(par_done_reg859_out),
      .done(par_done_reg859_done)
  );
  
  std_reg #(1) par_done_reg860 (
      .in(par_done_reg860_in),
      .write_en(par_done_reg860_write_en),
      .clk(clk),
      .out(par_done_reg860_out),
      .done(par_done_reg860_done)
  );
  
  std_reg #(1) par_done_reg861 (
      .in(par_done_reg861_in),
      .write_en(par_done_reg861_write_en),
      .clk(clk),
      .out(par_done_reg861_out),
      .done(par_done_reg861_done)
  );
  
  std_reg #(1) par_done_reg862 (
      .in(par_done_reg862_in),
      .write_en(par_done_reg862_write_en),
      .clk(clk),
      .out(par_done_reg862_out),
      .done(par_done_reg862_done)
  );
  
  std_reg #(1) par_done_reg863 (
      .in(par_done_reg863_in),
      .write_en(par_done_reg863_write_en),
      .clk(clk),
      .out(par_done_reg863_out),
      .done(par_done_reg863_done)
  );
  
  std_reg #(1) par_done_reg864 (
      .in(par_done_reg864_in),
      .write_en(par_done_reg864_write_en),
      .clk(clk),
      .out(par_done_reg864_out),
      .done(par_done_reg864_done)
  );
  
  std_reg #(1) par_done_reg865 (
      .in(par_done_reg865_in),
      .write_en(par_done_reg865_write_en),
      .clk(clk),
      .out(par_done_reg865_out),
      .done(par_done_reg865_done)
  );
  
  std_reg #(1) par_done_reg866 (
      .in(par_done_reg866_in),
      .write_en(par_done_reg866_write_en),
      .clk(clk),
      .out(par_done_reg866_out),
      .done(par_done_reg866_done)
  );
  
  std_reg #(1) par_done_reg867 (
      .in(par_done_reg867_in),
      .write_en(par_done_reg867_write_en),
      .clk(clk),
      .out(par_done_reg867_out),
      .done(par_done_reg867_done)
  );
  
  std_reg #(1) par_done_reg868 (
      .in(par_done_reg868_in),
      .write_en(par_done_reg868_write_en),
      .clk(clk),
      .out(par_done_reg868_out),
      .done(par_done_reg868_done)
  );
  
  std_reg #(1) par_done_reg869 (
      .in(par_done_reg869_in),
      .write_en(par_done_reg869_write_en),
      .clk(clk),
      .out(par_done_reg869_out),
      .done(par_done_reg869_done)
  );
  
  std_reg #(1) par_done_reg870 (
      .in(par_done_reg870_in),
      .write_en(par_done_reg870_write_en),
      .clk(clk),
      .out(par_done_reg870_out),
      .done(par_done_reg870_done)
  );
  
  std_reg #(1) par_done_reg871 (
      .in(par_done_reg871_in),
      .write_en(par_done_reg871_write_en),
      .clk(clk),
      .out(par_done_reg871_out),
      .done(par_done_reg871_done)
  );
  
  std_reg #(1) par_done_reg872 (
      .in(par_done_reg872_in),
      .write_en(par_done_reg872_write_en),
      .clk(clk),
      .out(par_done_reg872_out),
      .done(par_done_reg872_done)
  );
  
  std_reg #(1) par_done_reg873 (
      .in(par_done_reg873_in),
      .write_en(par_done_reg873_write_en),
      .clk(clk),
      .out(par_done_reg873_out),
      .done(par_done_reg873_done)
  );
  
  std_reg #(1) par_done_reg874 (
      .in(par_done_reg874_in),
      .write_en(par_done_reg874_write_en),
      .clk(clk),
      .out(par_done_reg874_out),
      .done(par_done_reg874_done)
  );
  
  std_reg #(1) par_done_reg875 (
      .in(par_done_reg875_in),
      .write_en(par_done_reg875_write_en),
      .clk(clk),
      .out(par_done_reg875_out),
      .done(par_done_reg875_done)
  );
  
  std_reg #(1) par_done_reg876 (
      .in(par_done_reg876_in),
      .write_en(par_done_reg876_write_en),
      .clk(clk),
      .out(par_done_reg876_out),
      .done(par_done_reg876_done)
  );
  
  std_reg #(1) par_done_reg877 (
      .in(par_done_reg877_in),
      .write_en(par_done_reg877_write_en),
      .clk(clk),
      .out(par_done_reg877_out),
      .done(par_done_reg877_done)
  );
  
  std_reg #(1) par_done_reg878 (
      .in(par_done_reg878_in),
      .write_en(par_done_reg878_write_en),
      .clk(clk),
      .out(par_done_reg878_out),
      .done(par_done_reg878_done)
  );
  
  std_reg #(1) par_done_reg879 (
      .in(par_done_reg879_in),
      .write_en(par_done_reg879_write_en),
      .clk(clk),
      .out(par_done_reg879_out),
      .done(par_done_reg879_done)
  );
  
  std_reg #(1) par_done_reg880 (
      .in(par_done_reg880_in),
      .write_en(par_done_reg880_write_en),
      .clk(clk),
      .out(par_done_reg880_out),
      .done(par_done_reg880_done)
  );
  
  std_reg #(1) par_done_reg881 (
      .in(par_done_reg881_in),
      .write_en(par_done_reg881_write_en),
      .clk(clk),
      .out(par_done_reg881_out),
      .done(par_done_reg881_done)
  );
  
  std_reg #(1) par_done_reg882 (
      .in(par_done_reg882_in),
      .write_en(par_done_reg882_write_en),
      .clk(clk),
      .out(par_done_reg882_out),
      .done(par_done_reg882_done)
  );
  
  std_reg #(1) par_done_reg883 (
      .in(par_done_reg883_in),
      .write_en(par_done_reg883_write_en),
      .clk(clk),
      .out(par_done_reg883_out),
      .done(par_done_reg883_done)
  );
  
  std_reg #(1) par_done_reg884 (
      .in(par_done_reg884_in),
      .write_en(par_done_reg884_write_en),
      .clk(clk),
      .out(par_done_reg884_out),
      .done(par_done_reg884_done)
  );
  
  std_reg #(1) par_done_reg885 (
      .in(par_done_reg885_in),
      .write_en(par_done_reg885_write_en),
      .clk(clk),
      .out(par_done_reg885_out),
      .done(par_done_reg885_done)
  );
  
  std_reg #(1) par_done_reg886 (
      .in(par_done_reg886_in),
      .write_en(par_done_reg886_write_en),
      .clk(clk),
      .out(par_done_reg886_out),
      .done(par_done_reg886_done)
  );
  
  std_reg #(1) par_done_reg887 (
      .in(par_done_reg887_in),
      .write_en(par_done_reg887_write_en),
      .clk(clk),
      .out(par_done_reg887_out),
      .done(par_done_reg887_done)
  );
  
  std_reg #(1) par_done_reg888 (
      .in(par_done_reg888_in),
      .write_en(par_done_reg888_write_en),
      .clk(clk),
      .out(par_done_reg888_out),
      .done(par_done_reg888_done)
  );
  
  std_reg #(1) par_done_reg889 (
      .in(par_done_reg889_in),
      .write_en(par_done_reg889_write_en),
      .clk(clk),
      .out(par_done_reg889_out),
      .done(par_done_reg889_done)
  );
  
  std_reg #(1) par_done_reg890 (
      .in(par_done_reg890_in),
      .write_en(par_done_reg890_write_en),
      .clk(clk),
      .out(par_done_reg890_out),
      .done(par_done_reg890_done)
  );
  
  std_reg #(1) par_done_reg891 (
      .in(par_done_reg891_in),
      .write_en(par_done_reg891_write_en),
      .clk(clk),
      .out(par_done_reg891_out),
      .done(par_done_reg891_done)
  );
  
  std_reg #(1) par_done_reg892 (
      .in(par_done_reg892_in),
      .write_en(par_done_reg892_write_en),
      .clk(clk),
      .out(par_done_reg892_out),
      .done(par_done_reg892_done)
  );
  
  std_reg #(1) par_done_reg893 (
      .in(par_done_reg893_in),
      .write_en(par_done_reg893_write_en),
      .clk(clk),
      .out(par_done_reg893_out),
      .done(par_done_reg893_done)
  );
  
  std_reg #(1) par_done_reg894 (
      .in(par_done_reg894_in),
      .write_en(par_done_reg894_write_en),
      .clk(clk),
      .out(par_done_reg894_out),
      .done(par_done_reg894_done)
  );
  
  std_reg #(1) par_done_reg895 (
      .in(par_done_reg895_in),
      .write_en(par_done_reg895_write_en),
      .clk(clk),
      .out(par_done_reg895_out),
      .done(par_done_reg895_done)
  );
  
  std_reg #(1) par_done_reg896 (
      .in(par_done_reg896_in),
      .write_en(par_done_reg896_write_en),
      .clk(clk),
      .out(par_done_reg896_out),
      .done(par_done_reg896_done)
  );
  
  std_reg #(1) par_done_reg897 (
      .in(par_done_reg897_in),
      .write_en(par_done_reg897_write_en),
      .clk(clk),
      .out(par_done_reg897_out),
      .done(par_done_reg897_done)
  );
  
  std_reg #(1) par_done_reg898 (
      .in(par_done_reg898_in),
      .write_en(par_done_reg898_write_en),
      .clk(clk),
      .out(par_done_reg898_out),
      .done(par_done_reg898_done)
  );
  
  std_reg #(1) par_done_reg899 (
      .in(par_done_reg899_in),
      .write_en(par_done_reg899_write_en),
      .clk(clk),
      .out(par_done_reg899_out),
      .done(par_done_reg899_done)
  );
  
  std_reg #(1) par_reset24 (
      .in(par_reset24_in),
      .write_en(par_reset24_write_en),
      .clk(clk),
      .out(par_reset24_out),
      .done(par_reset24_done)
  );
  
  std_reg #(1) par_done_reg900 (
      .in(par_done_reg900_in),
      .write_en(par_done_reg900_write_en),
      .clk(clk),
      .out(par_done_reg900_out),
      .done(par_done_reg900_done)
  );
  
  std_reg #(1) par_done_reg901 (
      .in(par_done_reg901_in),
      .write_en(par_done_reg901_write_en),
      .clk(clk),
      .out(par_done_reg901_out),
      .done(par_done_reg901_done)
  );
  
  std_reg #(1) par_done_reg902 (
      .in(par_done_reg902_in),
      .write_en(par_done_reg902_write_en),
      .clk(clk),
      .out(par_done_reg902_out),
      .done(par_done_reg902_done)
  );
  
  std_reg #(1) par_done_reg903 (
      .in(par_done_reg903_in),
      .write_en(par_done_reg903_write_en),
      .clk(clk),
      .out(par_done_reg903_out),
      .done(par_done_reg903_done)
  );
  
  std_reg #(1) par_done_reg904 (
      .in(par_done_reg904_in),
      .write_en(par_done_reg904_write_en),
      .clk(clk),
      .out(par_done_reg904_out),
      .done(par_done_reg904_done)
  );
  
  std_reg #(1) par_done_reg905 (
      .in(par_done_reg905_in),
      .write_en(par_done_reg905_write_en),
      .clk(clk),
      .out(par_done_reg905_out),
      .done(par_done_reg905_done)
  );
  
  std_reg #(1) par_done_reg906 (
      .in(par_done_reg906_in),
      .write_en(par_done_reg906_write_en),
      .clk(clk),
      .out(par_done_reg906_out),
      .done(par_done_reg906_done)
  );
  
  std_reg #(1) par_done_reg907 (
      .in(par_done_reg907_in),
      .write_en(par_done_reg907_write_en),
      .clk(clk),
      .out(par_done_reg907_out),
      .done(par_done_reg907_done)
  );
  
  std_reg #(1) par_done_reg908 (
      .in(par_done_reg908_in),
      .write_en(par_done_reg908_write_en),
      .clk(clk),
      .out(par_done_reg908_out),
      .done(par_done_reg908_done)
  );
  
  std_reg #(1) par_done_reg909 (
      .in(par_done_reg909_in),
      .write_en(par_done_reg909_write_en),
      .clk(clk),
      .out(par_done_reg909_out),
      .done(par_done_reg909_done)
  );
  
  std_reg #(1) par_done_reg910 (
      .in(par_done_reg910_in),
      .write_en(par_done_reg910_write_en),
      .clk(clk),
      .out(par_done_reg910_out),
      .done(par_done_reg910_done)
  );
  
  std_reg #(1) par_done_reg911 (
      .in(par_done_reg911_in),
      .write_en(par_done_reg911_write_en),
      .clk(clk),
      .out(par_done_reg911_out),
      .done(par_done_reg911_done)
  );
  
  std_reg #(1) par_done_reg912 (
      .in(par_done_reg912_in),
      .write_en(par_done_reg912_write_en),
      .clk(clk),
      .out(par_done_reg912_out),
      .done(par_done_reg912_done)
  );
  
  std_reg #(1) par_done_reg913 (
      .in(par_done_reg913_in),
      .write_en(par_done_reg913_write_en),
      .clk(clk),
      .out(par_done_reg913_out),
      .done(par_done_reg913_done)
  );
  
  std_reg #(1) par_done_reg914 (
      .in(par_done_reg914_in),
      .write_en(par_done_reg914_write_en),
      .clk(clk),
      .out(par_done_reg914_out),
      .done(par_done_reg914_done)
  );
  
  std_reg #(1) par_done_reg915 (
      .in(par_done_reg915_in),
      .write_en(par_done_reg915_write_en),
      .clk(clk),
      .out(par_done_reg915_out),
      .done(par_done_reg915_done)
  );
  
  std_reg #(1) par_done_reg916 (
      .in(par_done_reg916_in),
      .write_en(par_done_reg916_write_en),
      .clk(clk),
      .out(par_done_reg916_out),
      .done(par_done_reg916_done)
  );
  
  std_reg #(1) par_done_reg917 (
      .in(par_done_reg917_in),
      .write_en(par_done_reg917_write_en),
      .clk(clk),
      .out(par_done_reg917_out),
      .done(par_done_reg917_done)
  );
  
  std_reg #(1) par_done_reg918 (
      .in(par_done_reg918_in),
      .write_en(par_done_reg918_write_en),
      .clk(clk),
      .out(par_done_reg918_out),
      .done(par_done_reg918_done)
  );
  
  std_reg #(1) par_done_reg919 (
      .in(par_done_reg919_in),
      .write_en(par_done_reg919_write_en),
      .clk(clk),
      .out(par_done_reg919_out),
      .done(par_done_reg919_done)
  );
  
  std_reg #(1) par_done_reg920 (
      .in(par_done_reg920_in),
      .write_en(par_done_reg920_write_en),
      .clk(clk),
      .out(par_done_reg920_out),
      .done(par_done_reg920_done)
  );
  
  std_reg #(1) par_done_reg921 (
      .in(par_done_reg921_in),
      .write_en(par_done_reg921_write_en),
      .clk(clk),
      .out(par_done_reg921_out),
      .done(par_done_reg921_done)
  );
  
  std_reg #(1) par_done_reg922 (
      .in(par_done_reg922_in),
      .write_en(par_done_reg922_write_en),
      .clk(clk),
      .out(par_done_reg922_out),
      .done(par_done_reg922_done)
  );
  
  std_reg #(1) par_done_reg923 (
      .in(par_done_reg923_in),
      .write_en(par_done_reg923_write_en),
      .clk(clk),
      .out(par_done_reg923_out),
      .done(par_done_reg923_done)
  );
  
  std_reg #(1) par_done_reg924 (
      .in(par_done_reg924_in),
      .write_en(par_done_reg924_write_en),
      .clk(clk),
      .out(par_done_reg924_out),
      .done(par_done_reg924_done)
  );
  
  std_reg #(1) par_done_reg925 (
      .in(par_done_reg925_in),
      .write_en(par_done_reg925_write_en),
      .clk(clk),
      .out(par_done_reg925_out),
      .done(par_done_reg925_done)
  );
  
  std_reg #(1) par_done_reg926 (
      .in(par_done_reg926_in),
      .write_en(par_done_reg926_write_en),
      .clk(clk),
      .out(par_done_reg926_out),
      .done(par_done_reg926_done)
  );
  
  std_reg #(1) par_done_reg927 (
      .in(par_done_reg927_in),
      .write_en(par_done_reg927_write_en),
      .clk(clk),
      .out(par_done_reg927_out),
      .done(par_done_reg927_done)
  );
  
  std_reg #(1) par_done_reg928 (
      .in(par_done_reg928_in),
      .write_en(par_done_reg928_write_en),
      .clk(clk),
      .out(par_done_reg928_out),
      .done(par_done_reg928_done)
  );
  
  std_reg #(1) par_done_reg929 (
      .in(par_done_reg929_in),
      .write_en(par_done_reg929_write_en),
      .clk(clk),
      .out(par_done_reg929_out),
      .done(par_done_reg929_done)
  );
  
  std_reg #(1) par_done_reg930 (
      .in(par_done_reg930_in),
      .write_en(par_done_reg930_write_en),
      .clk(clk),
      .out(par_done_reg930_out),
      .done(par_done_reg930_done)
  );
  
  std_reg #(1) par_done_reg931 (
      .in(par_done_reg931_in),
      .write_en(par_done_reg931_write_en),
      .clk(clk),
      .out(par_done_reg931_out),
      .done(par_done_reg931_done)
  );
  
  std_reg #(1) par_done_reg932 (
      .in(par_done_reg932_in),
      .write_en(par_done_reg932_write_en),
      .clk(clk),
      .out(par_done_reg932_out),
      .done(par_done_reg932_done)
  );
  
  std_reg #(1) par_done_reg933 (
      .in(par_done_reg933_in),
      .write_en(par_done_reg933_write_en),
      .clk(clk),
      .out(par_done_reg933_out),
      .done(par_done_reg933_done)
  );
  
  std_reg #(1) par_done_reg934 (
      .in(par_done_reg934_in),
      .write_en(par_done_reg934_write_en),
      .clk(clk),
      .out(par_done_reg934_out),
      .done(par_done_reg934_done)
  );
  
  std_reg #(1) par_done_reg935 (
      .in(par_done_reg935_in),
      .write_en(par_done_reg935_write_en),
      .clk(clk),
      .out(par_done_reg935_out),
      .done(par_done_reg935_done)
  );
  
  std_reg #(1) par_done_reg936 (
      .in(par_done_reg936_in),
      .write_en(par_done_reg936_write_en),
      .clk(clk),
      .out(par_done_reg936_out),
      .done(par_done_reg936_done)
  );
  
  std_reg #(1) par_done_reg937 (
      .in(par_done_reg937_in),
      .write_en(par_done_reg937_write_en),
      .clk(clk),
      .out(par_done_reg937_out),
      .done(par_done_reg937_done)
  );
  
  std_reg #(1) par_done_reg938 (
      .in(par_done_reg938_in),
      .write_en(par_done_reg938_write_en),
      .clk(clk),
      .out(par_done_reg938_out),
      .done(par_done_reg938_done)
  );
  
  std_reg #(1) par_done_reg939 (
      .in(par_done_reg939_in),
      .write_en(par_done_reg939_write_en),
      .clk(clk),
      .out(par_done_reg939_out),
      .done(par_done_reg939_done)
  );
  
  std_reg #(1) par_done_reg940 (
      .in(par_done_reg940_in),
      .write_en(par_done_reg940_write_en),
      .clk(clk),
      .out(par_done_reg940_out),
      .done(par_done_reg940_done)
  );
  
  std_reg #(1) par_done_reg941 (
      .in(par_done_reg941_in),
      .write_en(par_done_reg941_write_en),
      .clk(clk),
      .out(par_done_reg941_out),
      .done(par_done_reg941_done)
  );
  
  std_reg #(1) par_done_reg942 (
      .in(par_done_reg942_in),
      .write_en(par_done_reg942_write_en),
      .clk(clk),
      .out(par_done_reg942_out),
      .done(par_done_reg942_done)
  );
  
  std_reg #(1) par_done_reg943 (
      .in(par_done_reg943_in),
      .write_en(par_done_reg943_write_en),
      .clk(clk),
      .out(par_done_reg943_out),
      .done(par_done_reg943_done)
  );
  
  std_reg #(1) par_done_reg944 (
      .in(par_done_reg944_in),
      .write_en(par_done_reg944_write_en),
      .clk(clk),
      .out(par_done_reg944_out),
      .done(par_done_reg944_done)
  );
  
  std_reg #(1) par_done_reg945 (
      .in(par_done_reg945_in),
      .write_en(par_done_reg945_write_en),
      .clk(clk),
      .out(par_done_reg945_out),
      .done(par_done_reg945_done)
  );
  
  std_reg #(1) par_done_reg946 (
      .in(par_done_reg946_in),
      .write_en(par_done_reg946_write_en),
      .clk(clk),
      .out(par_done_reg946_out),
      .done(par_done_reg946_done)
  );
  
  std_reg #(1) par_done_reg947 (
      .in(par_done_reg947_in),
      .write_en(par_done_reg947_write_en),
      .clk(clk),
      .out(par_done_reg947_out),
      .done(par_done_reg947_done)
  );
  
  std_reg #(1) par_done_reg948 (
      .in(par_done_reg948_in),
      .write_en(par_done_reg948_write_en),
      .clk(clk),
      .out(par_done_reg948_out),
      .done(par_done_reg948_done)
  );
  
  std_reg #(1) par_done_reg949 (
      .in(par_done_reg949_in),
      .write_en(par_done_reg949_write_en),
      .clk(clk),
      .out(par_done_reg949_out),
      .done(par_done_reg949_done)
  );
  
  std_reg #(1) par_done_reg950 (
      .in(par_done_reg950_in),
      .write_en(par_done_reg950_write_en),
      .clk(clk),
      .out(par_done_reg950_out),
      .done(par_done_reg950_done)
  );
  
  std_reg #(1) par_done_reg951 (
      .in(par_done_reg951_in),
      .write_en(par_done_reg951_write_en),
      .clk(clk),
      .out(par_done_reg951_out),
      .done(par_done_reg951_done)
  );
  
  std_reg #(1) par_done_reg952 (
      .in(par_done_reg952_in),
      .write_en(par_done_reg952_write_en),
      .clk(clk),
      .out(par_done_reg952_out),
      .done(par_done_reg952_done)
  );
  
  std_reg #(1) par_done_reg953 (
      .in(par_done_reg953_in),
      .write_en(par_done_reg953_write_en),
      .clk(clk),
      .out(par_done_reg953_out),
      .done(par_done_reg953_done)
  );
  
  std_reg #(1) par_done_reg954 (
      .in(par_done_reg954_in),
      .write_en(par_done_reg954_write_en),
      .clk(clk),
      .out(par_done_reg954_out),
      .done(par_done_reg954_done)
  );
  
  std_reg #(1) par_done_reg955 (
      .in(par_done_reg955_in),
      .write_en(par_done_reg955_write_en),
      .clk(clk),
      .out(par_done_reg955_out),
      .done(par_done_reg955_done)
  );
  
  std_reg #(1) par_done_reg956 (
      .in(par_done_reg956_in),
      .write_en(par_done_reg956_write_en),
      .clk(clk),
      .out(par_done_reg956_out),
      .done(par_done_reg956_done)
  );
  
  std_reg #(1) par_done_reg957 (
      .in(par_done_reg957_in),
      .write_en(par_done_reg957_write_en),
      .clk(clk),
      .out(par_done_reg957_out),
      .done(par_done_reg957_done)
  );
  
  std_reg #(1) par_done_reg958 (
      .in(par_done_reg958_in),
      .write_en(par_done_reg958_write_en),
      .clk(clk),
      .out(par_done_reg958_out),
      .done(par_done_reg958_done)
  );
  
  std_reg #(1) par_done_reg959 (
      .in(par_done_reg959_in),
      .write_en(par_done_reg959_write_en),
      .clk(clk),
      .out(par_done_reg959_out),
      .done(par_done_reg959_done)
  );
  
  std_reg #(1) par_done_reg960 (
      .in(par_done_reg960_in),
      .write_en(par_done_reg960_write_en),
      .clk(clk),
      .out(par_done_reg960_out),
      .done(par_done_reg960_done)
  );
  
  std_reg #(1) par_done_reg961 (
      .in(par_done_reg961_in),
      .write_en(par_done_reg961_write_en),
      .clk(clk),
      .out(par_done_reg961_out),
      .done(par_done_reg961_done)
  );
  
  std_reg #(1) par_done_reg962 (
      .in(par_done_reg962_in),
      .write_en(par_done_reg962_write_en),
      .clk(clk),
      .out(par_done_reg962_out),
      .done(par_done_reg962_done)
  );
  
  std_reg #(1) par_done_reg963 (
      .in(par_done_reg963_in),
      .write_en(par_done_reg963_write_en),
      .clk(clk),
      .out(par_done_reg963_out),
      .done(par_done_reg963_done)
  );
  
  std_reg #(1) par_done_reg964 (
      .in(par_done_reg964_in),
      .write_en(par_done_reg964_write_en),
      .clk(clk),
      .out(par_done_reg964_out),
      .done(par_done_reg964_done)
  );
  
  std_reg #(1) par_done_reg965 (
      .in(par_done_reg965_in),
      .write_en(par_done_reg965_write_en),
      .clk(clk),
      .out(par_done_reg965_out),
      .done(par_done_reg965_done)
  );
  
  std_reg #(1) par_done_reg966 (
      .in(par_done_reg966_in),
      .write_en(par_done_reg966_write_en),
      .clk(clk),
      .out(par_done_reg966_out),
      .done(par_done_reg966_done)
  );
  
  std_reg #(1) par_done_reg967 (
      .in(par_done_reg967_in),
      .write_en(par_done_reg967_write_en),
      .clk(clk),
      .out(par_done_reg967_out),
      .done(par_done_reg967_done)
  );
  
  std_reg #(1) par_done_reg968 (
      .in(par_done_reg968_in),
      .write_en(par_done_reg968_write_en),
      .clk(clk),
      .out(par_done_reg968_out),
      .done(par_done_reg968_done)
  );
  
  std_reg #(1) par_done_reg969 (
      .in(par_done_reg969_in),
      .write_en(par_done_reg969_write_en),
      .clk(clk),
      .out(par_done_reg969_out),
      .done(par_done_reg969_done)
  );
  
  std_reg #(1) par_done_reg970 (
      .in(par_done_reg970_in),
      .write_en(par_done_reg970_write_en),
      .clk(clk),
      .out(par_done_reg970_out),
      .done(par_done_reg970_done)
  );
  
  std_reg #(1) par_done_reg971 (
      .in(par_done_reg971_in),
      .write_en(par_done_reg971_write_en),
      .clk(clk),
      .out(par_done_reg971_out),
      .done(par_done_reg971_done)
  );
  
  std_reg #(1) par_done_reg972 (
      .in(par_done_reg972_in),
      .write_en(par_done_reg972_write_en),
      .clk(clk),
      .out(par_done_reg972_out),
      .done(par_done_reg972_done)
  );
  
  std_reg #(1) par_done_reg973 (
      .in(par_done_reg973_in),
      .write_en(par_done_reg973_write_en),
      .clk(clk),
      .out(par_done_reg973_out),
      .done(par_done_reg973_done)
  );
  
  std_reg #(1) par_done_reg974 (
      .in(par_done_reg974_in),
      .write_en(par_done_reg974_write_en),
      .clk(clk),
      .out(par_done_reg974_out),
      .done(par_done_reg974_done)
  );
  
  std_reg #(1) par_done_reg975 (
      .in(par_done_reg975_in),
      .write_en(par_done_reg975_write_en),
      .clk(clk),
      .out(par_done_reg975_out),
      .done(par_done_reg975_done)
  );
  
  std_reg #(1) par_done_reg976 (
      .in(par_done_reg976_in),
      .write_en(par_done_reg976_write_en),
      .clk(clk),
      .out(par_done_reg976_out),
      .done(par_done_reg976_done)
  );
  
  std_reg #(1) par_done_reg977 (
      .in(par_done_reg977_in),
      .write_en(par_done_reg977_write_en),
      .clk(clk),
      .out(par_done_reg977_out),
      .done(par_done_reg977_done)
  );
  
  std_reg #(1) par_done_reg978 (
      .in(par_done_reg978_in),
      .write_en(par_done_reg978_write_en),
      .clk(clk),
      .out(par_done_reg978_out),
      .done(par_done_reg978_done)
  );
  
  std_reg #(1) par_done_reg979 (
      .in(par_done_reg979_in),
      .write_en(par_done_reg979_write_en),
      .clk(clk),
      .out(par_done_reg979_out),
      .done(par_done_reg979_done)
  );
  
  std_reg #(1) par_done_reg980 (
      .in(par_done_reg980_in),
      .write_en(par_done_reg980_write_en),
      .clk(clk),
      .out(par_done_reg980_out),
      .done(par_done_reg980_done)
  );
  
  std_reg #(1) par_done_reg981 (
      .in(par_done_reg981_in),
      .write_en(par_done_reg981_write_en),
      .clk(clk),
      .out(par_done_reg981_out),
      .done(par_done_reg981_done)
  );
  
  std_reg #(1) par_done_reg982 (
      .in(par_done_reg982_in),
      .write_en(par_done_reg982_write_en),
      .clk(clk),
      .out(par_done_reg982_out),
      .done(par_done_reg982_done)
  );
  
  std_reg #(1) par_done_reg983 (
      .in(par_done_reg983_in),
      .write_en(par_done_reg983_write_en),
      .clk(clk),
      .out(par_done_reg983_out),
      .done(par_done_reg983_done)
  );
  
  std_reg #(1) par_done_reg984 (
      .in(par_done_reg984_in),
      .write_en(par_done_reg984_write_en),
      .clk(clk),
      .out(par_done_reg984_out),
      .done(par_done_reg984_done)
  );
  
  std_reg #(1) par_done_reg985 (
      .in(par_done_reg985_in),
      .write_en(par_done_reg985_write_en),
      .clk(clk),
      .out(par_done_reg985_out),
      .done(par_done_reg985_done)
  );
  
  std_reg #(1) par_done_reg986 (
      .in(par_done_reg986_in),
      .write_en(par_done_reg986_write_en),
      .clk(clk),
      .out(par_done_reg986_out),
      .done(par_done_reg986_done)
  );
  
  std_reg #(1) par_done_reg987 (
      .in(par_done_reg987_in),
      .write_en(par_done_reg987_write_en),
      .clk(clk),
      .out(par_done_reg987_out),
      .done(par_done_reg987_done)
  );
  
  std_reg #(1) par_done_reg988 (
      .in(par_done_reg988_in),
      .write_en(par_done_reg988_write_en),
      .clk(clk),
      .out(par_done_reg988_out),
      .done(par_done_reg988_done)
  );
  
  std_reg #(1) par_done_reg989 (
      .in(par_done_reg989_in),
      .write_en(par_done_reg989_write_en),
      .clk(clk),
      .out(par_done_reg989_out),
      .done(par_done_reg989_done)
  );
  
  std_reg #(1) par_done_reg990 (
      .in(par_done_reg990_in),
      .write_en(par_done_reg990_write_en),
      .clk(clk),
      .out(par_done_reg990_out),
      .done(par_done_reg990_done)
  );
  
  std_reg #(1) par_done_reg991 (
      .in(par_done_reg991_in),
      .write_en(par_done_reg991_write_en),
      .clk(clk),
      .out(par_done_reg991_out),
      .done(par_done_reg991_done)
  );
  
  std_reg #(1) par_done_reg992 (
      .in(par_done_reg992_in),
      .write_en(par_done_reg992_write_en),
      .clk(clk),
      .out(par_done_reg992_out),
      .done(par_done_reg992_done)
  );
  
  std_reg #(1) par_done_reg993 (
      .in(par_done_reg993_in),
      .write_en(par_done_reg993_write_en),
      .clk(clk),
      .out(par_done_reg993_out),
      .done(par_done_reg993_done)
  );
  
  std_reg #(1) par_done_reg994 (
      .in(par_done_reg994_in),
      .write_en(par_done_reg994_write_en),
      .clk(clk),
      .out(par_done_reg994_out),
      .done(par_done_reg994_done)
  );
  
  std_reg #(1) par_done_reg995 (
      .in(par_done_reg995_in),
      .write_en(par_done_reg995_write_en),
      .clk(clk),
      .out(par_done_reg995_out),
      .done(par_done_reg995_done)
  );
  
  std_reg #(1) par_reset25 (
      .in(par_reset25_in),
      .write_en(par_reset25_write_en),
      .clk(clk),
      .out(par_reset25_out),
      .done(par_reset25_done)
  );
  
  std_reg #(1) par_done_reg996 (
      .in(par_done_reg996_in),
      .write_en(par_done_reg996_write_en),
      .clk(clk),
      .out(par_done_reg996_out),
      .done(par_done_reg996_done)
  );
  
  std_reg #(1) par_done_reg997 (
      .in(par_done_reg997_in),
      .write_en(par_done_reg997_write_en),
      .clk(clk),
      .out(par_done_reg997_out),
      .done(par_done_reg997_done)
  );
  
  std_reg #(1) par_done_reg998 (
      .in(par_done_reg998_in),
      .write_en(par_done_reg998_write_en),
      .clk(clk),
      .out(par_done_reg998_out),
      .done(par_done_reg998_done)
  );
  
  std_reg #(1) par_done_reg999 (
      .in(par_done_reg999_in),
      .write_en(par_done_reg999_write_en),
      .clk(clk),
      .out(par_done_reg999_out),
      .done(par_done_reg999_done)
  );
  
  std_reg #(1) par_done_reg1000 (
      .in(par_done_reg1000_in),
      .write_en(par_done_reg1000_write_en),
      .clk(clk),
      .out(par_done_reg1000_out),
      .done(par_done_reg1000_done)
  );
  
  std_reg #(1) par_done_reg1001 (
      .in(par_done_reg1001_in),
      .write_en(par_done_reg1001_write_en),
      .clk(clk),
      .out(par_done_reg1001_out),
      .done(par_done_reg1001_done)
  );
  
  std_reg #(1) par_done_reg1002 (
      .in(par_done_reg1002_in),
      .write_en(par_done_reg1002_write_en),
      .clk(clk),
      .out(par_done_reg1002_out),
      .done(par_done_reg1002_done)
  );
  
  std_reg #(1) par_done_reg1003 (
      .in(par_done_reg1003_in),
      .write_en(par_done_reg1003_write_en),
      .clk(clk),
      .out(par_done_reg1003_out),
      .done(par_done_reg1003_done)
  );
  
  std_reg #(1) par_done_reg1004 (
      .in(par_done_reg1004_in),
      .write_en(par_done_reg1004_write_en),
      .clk(clk),
      .out(par_done_reg1004_out),
      .done(par_done_reg1004_done)
  );
  
  std_reg #(1) par_done_reg1005 (
      .in(par_done_reg1005_in),
      .write_en(par_done_reg1005_write_en),
      .clk(clk),
      .out(par_done_reg1005_out),
      .done(par_done_reg1005_done)
  );
  
  std_reg #(1) par_done_reg1006 (
      .in(par_done_reg1006_in),
      .write_en(par_done_reg1006_write_en),
      .clk(clk),
      .out(par_done_reg1006_out),
      .done(par_done_reg1006_done)
  );
  
  std_reg #(1) par_done_reg1007 (
      .in(par_done_reg1007_in),
      .write_en(par_done_reg1007_write_en),
      .clk(clk),
      .out(par_done_reg1007_out),
      .done(par_done_reg1007_done)
  );
  
  std_reg #(1) par_done_reg1008 (
      .in(par_done_reg1008_in),
      .write_en(par_done_reg1008_write_en),
      .clk(clk),
      .out(par_done_reg1008_out),
      .done(par_done_reg1008_done)
  );
  
  std_reg #(1) par_done_reg1009 (
      .in(par_done_reg1009_in),
      .write_en(par_done_reg1009_write_en),
      .clk(clk),
      .out(par_done_reg1009_out),
      .done(par_done_reg1009_done)
  );
  
  std_reg #(1) par_done_reg1010 (
      .in(par_done_reg1010_in),
      .write_en(par_done_reg1010_write_en),
      .clk(clk),
      .out(par_done_reg1010_out),
      .done(par_done_reg1010_done)
  );
  
  std_reg #(1) par_done_reg1011 (
      .in(par_done_reg1011_in),
      .write_en(par_done_reg1011_write_en),
      .clk(clk),
      .out(par_done_reg1011_out),
      .done(par_done_reg1011_done)
  );
  
  std_reg #(1) par_done_reg1012 (
      .in(par_done_reg1012_in),
      .write_en(par_done_reg1012_write_en),
      .clk(clk),
      .out(par_done_reg1012_out),
      .done(par_done_reg1012_done)
  );
  
  std_reg #(1) par_done_reg1013 (
      .in(par_done_reg1013_in),
      .write_en(par_done_reg1013_write_en),
      .clk(clk),
      .out(par_done_reg1013_out),
      .done(par_done_reg1013_done)
  );
  
  std_reg #(1) par_done_reg1014 (
      .in(par_done_reg1014_in),
      .write_en(par_done_reg1014_write_en),
      .clk(clk),
      .out(par_done_reg1014_out),
      .done(par_done_reg1014_done)
  );
  
  std_reg #(1) par_done_reg1015 (
      .in(par_done_reg1015_in),
      .write_en(par_done_reg1015_write_en),
      .clk(clk),
      .out(par_done_reg1015_out),
      .done(par_done_reg1015_done)
  );
  
  std_reg #(1) par_done_reg1016 (
      .in(par_done_reg1016_in),
      .write_en(par_done_reg1016_write_en),
      .clk(clk),
      .out(par_done_reg1016_out),
      .done(par_done_reg1016_done)
  );
  
  std_reg #(1) par_done_reg1017 (
      .in(par_done_reg1017_in),
      .write_en(par_done_reg1017_write_en),
      .clk(clk),
      .out(par_done_reg1017_out),
      .done(par_done_reg1017_done)
  );
  
  std_reg #(1) par_done_reg1018 (
      .in(par_done_reg1018_in),
      .write_en(par_done_reg1018_write_en),
      .clk(clk),
      .out(par_done_reg1018_out),
      .done(par_done_reg1018_done)
  );
  
  std_reg #(1) par_done_reg1019 (
      .in(par_done_reg1019_in),
      .write_en(par_done_reg1019_write_en),
      .clk(clk),
      .out(par_done_reg1019_out),
      .done(par_done_reg1019_done)
  );
  
  std_reg #(1) par_done_reg1020 (
      .in(par_done_reg1020_in),
      .write_en(par_done_reg1020_write_en),
      .clk(clk),
      .out(par_done_reg1020_out),
      .done(par_done_reg1020_done)
  );
  
  std_reg #(1) par_done_reg1021 (
      .in(par_done_reg1021_in),
      .write_en(par_done_reg1021_write_en),
      .clk(clk),
      .out(par_done_reg1021_out),
      .done(par_done_reg1021_done)
  );
  
  std_reg #(1) par_done_reg1022 (
      .in(par_done_reg1022_in),
      .write_en(par_done_reg1022_write_en),
      .clk(clk),
      .out(par_done_reg1022_out),
      .done(par_done_reg1022_done)
  );
  
  std_reg #(1) par_done_reg1023 (
      .in(par_done_reg1023_in),
      .write_en(par_done_reg1023_write_en),
      .clk(clk),
      .out(par_done_reg1023_out),
      .done(par_done_reg1023_done)
  );
  
  std_reg #(1) par_done_reg1024 (
      .in(par_done_reg1024_in),
      .write_en(par_done_reg1024_write_en),
      .clk(clk),
      .out(par_done_reg1024_out),
      .done(par_done_reg1024_done)
  );
  
  std_reg #(1) par_done_reg1025 (
      .in(par_done_reg1025_in),
      .write_en(par_done_reg1025_write_en),
      .clk(clk),
      .out(par_done_reg1025_out),
      .done(par_done_reg1025_done)
  );
  
  std_reg #(1) par_done_reg1026 (
      .in(par_done_reg1026_in),
      .write_en(par_done_reg1026_write_en),
      .clk(clk),
      .out(par_done_reg1026_out),
      .done(par_done_reg1026_done)
  );
  
  std_reg #(1) par_done_reg1027 (
      .in(par_done_reg1027_in),
      .write_en(par_done_reg1027_write_en),
      .clk(clk),
      .out(par_done_reg1027_out),
      .done(par_done_reg1027_done)
  );
  
  std_reg #(1) par_done_reg1028 (
      .in(par_done_reg1028_in),
      .write_en(par_done_reg1028_write_en),
      .clk(clk),
      .out(par_done_reg1028_out),
      .done(par_done_reg1028_done)
  );
  
  std_reg #(1) par_done_reg1029 (
      .in(par_done_reg1029_in),
      .write_en(par_done_reg1029_write_en),
      .clk(clk),
      .out(par_done_reg1029_out),
      .done(par_done_reg1029_done)
  );
  
  std_reg #(1) par_done_reg1030 (
      .in(par_done_reg1030_in),
      .write_en(par_done_reg1030_write_en),
      .clk(clk),
      .out(par_done_reg1030_out),
      .done(par_done_reg1030_done)
  );
  
  std_reg #(1) par_done_reg1031 (
      .in(par_done_reg1031_in),
      .write_en(par_done_reg1031_write_en),
      .clk(clk),
      .out(par_done_reg1031_out),
      .done(par_done_reg1031_done)
  );
  
  std_reg #(1) par_done_reg1032 (
      .in(par_done_reg1032_in),
      .write_en(par_done_reg1032_write_en),
      .clk(clk),
      .out(par_done_reg1032_out),
      .done(par_done_reg1032_done)
  );
  
  std_reg #(1) par_done_reg1033 (
      .in(par_done_reg1033_in),
      .write_en(par_done_reg1033_write_en),
      .clk(clk),
      .out(par_done_reg1033_out),
      .done(par_done_reg1033_done)
  );
  
  std_reg #(1) par_done_reg1034 (
      .in(par_done_reg1034_in),
      .write_en(par_done_reg1034_write_en),
      .clk(clk),
      .out(par_done_reg1034_out),
      .done(par_done_reg1034_done)
  );
  
  std_reg #(1) par_done_reg1035 (
      .in(par_done_reg1035_in),
      .write_en(par_done_reg1035_write_en),
      .clk(clk),
      .out(par_done_reg1035_out),
      .done(par_done_reg1035_done)
  );
  
  std_reg #(1) par_done_reg1036 (
      .in(par_done_reg1036_in),
      .write_en(par_done_reg1036_write_en),
      .clk(clk),
      .out(par_done_reg1036_out),
      .done(par_done_reg1036_done)
  );
  
  std_reg #(1) par_done_reg1037 (
      .in(par_done_reg1037_in),
      .write_en(par_done_reg1037_write_en),
      .clk(clk),
      .out(par_done_reg1037_out),
      .done(par_done_reg1037_done)
  );
  
  std_reg #(1) par_done_reg1038 (
      .in(par_done_reg1038_in),
      .write_en(par_done_reg1038_write_en),
      .clk(clk),
      .out(par_done_reg1038_out),
      .done(par_done_reg1038_done)
  );
  
  std_reg #(1) par_done_reg1039 (
      .in(par_done_reg1039_in),
      .write_en(par_done_reg1039_write_en),
      .clk(clk),
      .out(par_done_reg1039_out),
      .done(par_done_reg1039_done)
  );
  
  std_reg #(1) par_done_reg1040 (
      .in(par_done_reg1040_in),
      .write_en(par_done_reg1040_write_en),
      .clk(clk),
      .out(par_done_reg1040_out),
      .done(par_done_reg1040_done)
  );
  
  std_reg #(1) par_done_reg1041 (
      .in(par_done_reg1041_in),
      .write_en(par_done_reg1041_write_en),
      .clk(clk),
      .out(par_done_reg1041_out),
      .done(par_done_reg1041_done)
  );
  
  std_reg #(1) par_done_reg1042 (
      .in(par_done_reg1042_in),
      .write_en(par_done_reg1042_write_en),
      .clk(clk),
      .out(par_done_reg1042_out),
      .done(par_done_reg1042_done)
  );
  
  std_reg #(1) par_done_reg1043 (
      .in(par_done_reg1043_in),
      .write_en(par_done_reg1043_write_en),
      .clk(clk),
      .out(par_done_reg1043_out),
      .done(par_done_reg1043_done)
  );
  
  std_reg #(1) par_done_reg1044 (
      .in(par_done_reg1044_in),
      .write_en(par_done_reg1044_write_en),
      .clk(clk),
      .out(par_done_reg1044_out),
      .done(par_done_reg1044_done)
  );
  
  std_reg #(1) par_done_reg1045 (
      .in(par_done_reg1045_in),
      .write_en(par_done_reg1045_write_en),
      .clk(clk),
      .out(par_done_reg1045_out),
      .done(par_done_reg1045_done)
  );
  
  std_reg #(1) par_done_reg1046 (
      .in(par_done_reg1046_in),
      .write_en(par_done_reg1046_write_en),
      .clk(clk),
      .out(par_done_reg1046_out),
      .done(par_done_reg1046_done)
  );
  
  std_reg #(1) par_done_reg1047 (
      .in(par_done_reg1047_in),
      .write_en(par_done_reg1047_write_en),
      .clk(clk),
      .out(par_done_reg1047_out),
      .done(par_done_reg1047_done)
  );
  
  std_reg #(1) par_done_reg1048 (
      .in(par_done_reg1048_in),
      .write_en(par_done_reg1048_write_en),
      .clk(clk),
      .out(par_done_reg1048_out),
      .done(par_done_reg1048_done)
  );
  
  std_reg #(1) par_done_reg1049 (
      .in(par_done_reg1049_in),
      .write_en(par_done_reg1049_write_en),
      .clk(clk),
      .out(par_done_reg1049_out),
      .done(par_done_reg1049_done)
  );
  
  std_reg #(1) par_reset26 (
      .in(par_reset26_in),
      .write_en(par_reset26_write_en),
      .clk(clk),
      .out(par_reset26_out),
      .done(par_reset26_done)
  );
  
  std_reg #(1) par_done_reg1050 (
      .in(par_done_reg1050_in),
      .write_en(par_done_reg1050_write_en),
      .clk(clk),
      .out(par_done_reg1050_out),
      .done(par_done_reg1050_done)
  );
  
  std_reg #(1) par_done_reg1051 (
      .in(par_done_reg1051_in),
      .write_en(par_done_reg1051_write_en),
      .clk(clk),
      .out(par_done_reg1051_out),
      .done(par_done_reg1051_done)
  );
  
  std_reg #(1) par_done_reg1052 (
      .in(par_done_reg1052_in),
      .write_en(par_done_reg1052_write_en),
      .clk(clk),
      .out(par_done_reg1052_out),
      .done(par_done_reg1052_done)
  );
  
  std_reg #(1) par_done_reg1053 (
      .in(par_done_reg1053_in),
      .write_en(par_done_reg1053_write_en),
      .clk(clk),
      .out(par_done_reg1053_out),
      .done(par_done_reg1053_done)
  );
  
  std_reg #(1) par_done_reg1054 (
      .in(par_done_reg1054_in),
      .write_en(par_done_reg1054_write_en),
      .clk(clk),
      .out(par_done_reg1054_out),
      .done(par_done_reg1054_done)
  );
  
  std_reg #(1) par_done_reg1055 (
      .in(par_done_reg1055_in),
      .write_en(par_done_reg1055_write_en),
      .clk(clk),
      .out(par_done_reg1055_out),
      .done(par_done_reg1055_done)
  );
  
  std_reg #(1) par_done_reg1056 (
      .in(par_done_reg1056_in),
      .write_en(par_done_reg1056_write_en),
      .clk(clk),
      .out(par_done_reg1056_out),
      .done(par_done_reg1056_done)
  );
  
  std_reg #(1) par_done_reg1057 (
      .in(par_done_reg1057_in),
      .write_en(par_done_reg1057_write_en),
      .clk(clk),
      .out(par_done_reg1057_out),
      .done(par_done_reg1057_done)
  );
  
  std_reg #(1) par_done_reg1058 (
      .in(par_done_reg1058_in),
      .write_en(par_done_reg1058_write_en),
      .clk(clk),
      .out(par_done_reg1058_out),
      .done(par_done_reg1058_done)
  );
  
  std_reg #(1) par_done_reg1059 (
      .in(par_done_reg1059_in),
      .write_en(par_done_reg1059_write_en),
      .clk(clk),
      .out(par_done_reg1059_out),
      .done(par_done_reg1059_done)
  );
  
  std_reg #(1) par_done_reg1060 (
      .in(par_done_reg1060_in),
      .write_en(par_done_reg1060_write_en),
      .clk(clk),
      .out(par_done_reg1060_out),
      .done(par_done_reg1060_done)
  );
  
  std_reg #(1) par_done_reg1061 (
      .in(par_done_reg1061_in),
      .write_en(par_done_reg1061_write_en),
      .clk(clk),
      .out(par_done_reg1061_out),
      .done(par_done_reg1061_done)
  );
  
  std_reg #(1) par_done_reg1062 (
      .in(par_done_reg1062_in),
      .write_en(par_done_reg1062_write_en),
      .clk(clk),
      .out(par_done_reg1062_out),
      .done(par_done_reg1062_done)
  );
  
  std_reg #(1) par_done_reg1063 (
      .in(par_done_reg1063_in),
      .write_en(par_done_reg1063_write_en),
      .clk(clk),
      .out(par_done_reg1063_out),
      .done(par_done_reg1063_done)
  );
  
  std_reg #(1) par_done_reg1064 (
      .in(par_done_reg1064_in),
      .write_en(par_done_reg1064_write_en),
      .clk(clk),
      .out(par_done_reg1064_out),
      .done(par_done_reg1064_done)
  );
  
  std_reg #(1) par_done_reg1065 (
      .in(par_done_reg1065_in),
      .write_en(par_done_reg1065_write_en),
      .clk(clk),
      .out(par_done_reg1065_out),
      .done(par_done_reg1065_done)
  );
  
  std_reg #(1) par_done_reg1066 (
      .in(par_done_reg1066_in),
      .write_en(par_done_reg1066_write_en),
      .clk(clk),
      .out(par_done_reg1066_out),
      .done(par_done_reg1066_done)
  );
  
  std_reg #(1) par_done_reg1067 (
      .in(par_done_reg1067_in),
      .write_en(par_done_reg1067_write_en),
      .clk(clk),
      .out(par_done_reg1067_out),
      .done(par_done_reg1067_done)
  );
  
  std_reg #(1) par_done_reg1068 (
      .in(par_done_reg1068_in),
      .write_en(par_done_reg1068_write_en),
      .clk(clk),
      .out(par_done_reg1068_out),
      .done(par_done_reg1068_done)
  );
  
  std_reg #(1) par_done_reg1069 (
      .in(par_done_reg1069_in),
      .write_en(par_done_reg1069_write_en),
      .clk(clk),
      .out(par_done_reg1069_out),
      .done(par_done_reg1069_done)
  );
  
  std_reg #(1) par_done_reg1070 (
      .in(par_done_reg1070_in),
      .write_en(par_done_reg1070_write_en),
      .clk(clk),
      .out(par_done_reg1070_out),
      .done(par_done_reg1070_done)
  );
  
  std_reg #(1) par_done_reg1071 (
      .in(par_done_reg1071_in),
      .write_en(par_done_reg1071_write_en),
      .clk(clk),
      .out(par_done_reg1071_out),
      .done(par_done_reg1071_done)
  );
  
  std_reg #(1) par_done_reg1072 (
      .in(par_done_reg1072_in),
      .write_en(par_done_reg1072_write_en),
      .clk(clk),
      .out(par_done_reg1072_out),
      .done(par_done_reg1072_done)
  );
  
  std_reg #(1) par_done_reg1073 (
      .in(par_done_reg1073_in),
      .write_en(par_done_reg1073_write_en),
      .clk(clk),
      .out(par_done_reg1073_out),
      .done(par_done_reg1073_done)
  );
  
  std_reg #(1) par_done_reg1074 (
      .in(par_done_reg1074_in),
      .write_en(par_done_reg1074_write_en),
      .clk(clk),
      .out(par_done_reg1074_out),
      .done(par_done_reg1074_done)
  );
  
  std_reg #(1) par_done_reg1075 (
      .in(par_done_reg1075_in),
      .write_en(par_done_reg1075_write_en),
      .clk(clk),
      .out(par_done_reg1075_out),
      .done(par_done_reg1075_done)
  );
  
  std_reg #(1) par_done_reg1076 (
      .in(par_done_reg1076_in),
      .write_en(par_done_reg1076_write_en),
      .clk(clk),
      .out(par_done_reg1076_out),
      .done(par_done_reg1076_done)
  );
  
  std_reg #(1) par_done_reg1077 (
      .in(par_done_reg1077_in),
      .write_en(par_done_reg1077_write_en),
      .clk(clk),
      .out(par_done_reg1077_out),
      .done(par_done_reg1077_done)
  );
  
  std_reg #(1) par_done_reg1078 (
      .in(par_done_reg1078_in),
      .write_en(par_done_reg1078_write_en),
      .clk(clk),
      .out(par_done_reg1078_out),
      .done(par_done_reg1078_done)
  );
  
  std_reg #(1) par_done_reg1079 (
      .in(par_done_reg1079_in),
      .write_en(par_done_reg1079_write_en),
      .clk(clk),
      .out(par_done_reg1079_out),
      .done(par_done_reg1079_done)
  );
  
  std_reg #(1) par_done_reg1080 (
      .in(par_done_reg1080_in),
      .write_en(par_done_reg1080_write_en),
      .clk(clk),
      .out(par_done_reg1080_out),
      .done(par_done_reg1080_done)
  );
  
  std_reg #(1) par_done_reg1081 (
      .in(par_done_reg1081_in),
      .write_en(par_done_reg1081_write_en),
      .clk(clk),
      .out(par_done_reg1081_out),
      .done(par_done_reg1081_done)
  );
  
  std_reg #(1) par_done_reg1082 (
      .in(par_done_reg1082_in),
      .write_en(par_done_reg1082_write_en),
      .clk(clk),
      .out(par_done_reg1082_out),
      .done(par_done_reg1082_done)
  );
  
  std_reg #(1) par_done_reg1083 (
      .in(par_done_reg1083_in),
      .write_en(par_done_reg1083_write_en),
      .clk(clk),
      .out(par_done_reg1083_out),
      .done(par_done_reg1083_done)
  );
  
  std_reg #(1) par_done_reg1084 (
      .in(par_done_reg1084_in),
      .write_en(par_done_reg1084_write_en),
      .clk(clk),
      .out(par_done_reg1084_out),
      .done(par_done_reg1084_done)
  );
  
  std_reg #(1) par_done_reg1085 (
      .in(par_done_reg1085_in),
      .write_en(par_done_reg1085_write_en),
      .clk(clk),
      .out(par_done_reg1085_out),
      .done(par_done_reg1085_done)
  );
  
  std_reg #(1) par_done_reg1086 (
      .in(par_done_reg1086_in),
      .write_en(par_done_reg1086_write_en),
      .clk(clk),
      .out(par_done_reg1086_out),
      .done(par_done_reg1086_done)
  );
  
  std_reg #(1) par_done_reg1087 (
      .in(par_done_reg1087_in),
      .write_en(par_done_reg1087_write_en),
      .clk(clk),
      .out(par_done_reg1087_out),
      .done(par_done_reg1087_done)
  );
  
  std_reg #(1) par_done_reg1088 (
      .in(par_done_reg1088_in),
      .write_en(par_done_reg1088_write_en),
      .clk(clk),
      .out(par_done_reg1088_out),
      .done(par_done_reg1088_done)
  );
  
  std_reg #(1) par_done_reg1089 (
      .in(par_done_reg1089_in),
      .write_en(par_done_reg1089_write_en),
      .clk(clk),
      .out(par_done_reg1089_out),
      .done(par_done_reg1089_done)
  );
  
  std_reg #(1) par_done_reg1090 (
      .in(par_done_reg1090_in),
      .write_en(par_done_reg1090_write_en),
      .clk(clk),
      .out(par_done_reg1090_out),
      .done(par_done_reg1090_done)
  );
  
  std_reg #(1) par_done_reg1091 (
      .in(par_done_reg1091_in),
      .write_en(par_done_reg1091_write_en),
      .clk(clk),
      .out(par_done_reg1091_out),
      .done(par_done_reg1091_done)
  );
  
  std_reg #(1) par_done_reg1092 (
      .in(par_done_reg1092_in),
      .write_en(par_done_reg1092_write_en),
      .clk(clk),
      .out(par_done_reg1092_out),
      .done(par_done_reg1092_done)
  );
  
  std_reg #(1) par_done_reg1093 (
      .in(par_done_reg1093_in),
      .write_en(par_done_reg1093_write_en),
      .clk(clk),
      .out(par_done_reg1093_out),
      .done(par_done_reg1093_done)
  );
  
  std_reg #(1) par_done_reg1094 (
      .in(par_done_reg1094_in),
      .write_en(par_done_reg1094_write_en),
      .clk(clk),
      .out(par_done_reg1094_out),
      .done(par_done_reg1094_done)
  );
  
  std_reg #(1) par_done_reg1095 (
      .in(par_done_reg1095_in),
      .write_en(par_done_reg1095_write_en),
      .clk(clk),
      .out(par_done_reg1095_out),
      .done(par_done_reg1095_done)
  );
  
  std_reg #(1) par_done_reg1096 (
      .in(par_done_reg1096_in),
      .write_en(par_done_reg1096_write_en),
      .clk(clk),
      .out(par_done_reg1096_out),
      .done(par_done_reg1096_done)
  );
  
  std_reg #(1) par_done_reg1097 (
      .in(par_done_reg1097_in),
      .write_en(par_done_reg1097_write_en),
      .clk(clk),
      .out(par_done_reg1097_out),
      .done(par_done_reg1097_done)
  );
  
  std_reg #(1) par_done_reg1098 (
      .in(par_done_reg1098_in),
      .write_en(par_done_reg1098_write_en),
      .clk(clk),
      .out(par_done_reg1098_out),
      .done(par_done_reg1098_done)
  );
  
  std_reg #(1) par_done_reg1099 (
      .in(par_done_reg1099_in),
      .write_en(par_done_reg1099_write_en),
      .clk(clk),
      .out(par_done_reg1099_out),
      .done(par_done_reg1099_done)
  );
  
  std_reg #(1) par_done_reg1100 (
      .in(par_done_reg1100_in),
      .write_en(par_done_reg1100_write_en),
      .clk(clk),
      .out(par_done_reg1100_out),
      .done(par_done_reg1100_done)
  );
  
  std_reg #(1) par_done_reg1101 (
      .in(par_done_reg1101_in),
      .write_en(par_done_reg1101_write_en),
      .clk(clk),
      .out(par_done_reg1101_out),
      .done(par_done_reg1101_done)
  );
  
  std_reg #(1) par_done_reg1102 (
      .in(par_done_reg1102_in),
      .write_en(par_done_reg1102_write_en),
      .clk(clk),
      .out(par_done_reg1102_out),
      .done(par_done_reg1102_done)
  );
  
  std_reg #(1) par_done_reg1103 (
      .in(par_done_reg1103_in),
      .write_en(par_done_reg1103_write_en),
      .clk(clk),
      .out(par_done_reg1103_out),
      .done(par_done_reg1103_done)
  );
  
  std_reg #(1) par_done_reg1104 (
      .in(par_done_reg1104_in),
      .write_en(par_done_reg1104_write_en),
      .clk(clk),
      .out(par_done_reg1104_out),
      .done(par_done_reg1104_done)
  );
  
  std_reg #(1) par_done_reg1105 (
      .in(par_done_reg1105_in),
      .write_en(par_done_reg1105_write_en),
      .clk(clk),
      .out(par_done_reg1105_out),
      .done(par_done_reg1105_done)
  );
  
  std_reg #(1) par_done_reg1106 (
      .in(par_done_reg1106_in),
      .write_en(par_done_reg1106_write_en),
      .clk(clk),
      .out(par_done_reg1106_out),
      .done(par_done_reg1106_done)
  );
  
  std_reg #(1) par_done_reg1107 (
      .in(par_done_reg1107_in),
      .write_en(par_done_reg1107_write_en),
      .clk(clk),
      .out(par_done_reg1107_out),
      .done(par_done_reg1107_done)
  );
  
  std_reg #(1) par_done_reg1108 (
      .in(par_done_reg1108_in),
      .write_en(par_done_reg1108_write_en),
      .clk(clk),
      .out(par_done_reg1108_out),
      .done(par_done_reg1108_done)
  );
  
  std_reg #(1) par_done_reg1109 (
      .in(par_done_reg1109_in),
      .write_en(par_done_reg1109_write_en),
      .clk(clk),
      .out(par_done_reg1109_out),
      .done(par_done_reg1109_done)
  );
  
  std_reg #(1) par_done_reg1110 (
      .in(par_done_reg1110_in),
      .write_en(par_done_reg1110_write_en),
      .clk(clk),
      .out(par_done_reg1110_out),
      .done(par_done_reg1110_done)
  );
  
  std_reg #(1) par_done_reg1111 (
      .in(par_done_reg1111_in),
      .write_en(par_done_reg1111_write_en),
      .clk(clk),
      .out(par_done_reg1111_out),
      .done(par_done_reg1111_done)
  );
  
  std_reg #(1) par_done_reg1112 (
      .in(par_done_reg1112_in),
      .write_en(par_done_reg1112_write_en),
      .clk(clk),
      .out(par_done_reg1112_out),
      .done(par_done_reg1112_done)
  );
  
  std_reg #(1) par_done_reg1113 (
      .in(par_done_reg1113_in),
      .write_en(par_done_reg1113_write_en),
      .clk(clk),
      .out(par_done_reg1113_out),
      .done(par_done_reg1113_done)
  );
  
  std_reg #(1) par_done_reg1114 (
      .in(par_done_reg1114_in),
      .write_en(par_done_reg1114_write_en),
      .clk(clk),
      .out(par_done_reg1114_out),
      .done(par_done_reg1114_done)
  );
  
  std_reg #(1) par_done_reg1115 (
      .in(par_done_reg1115_in),
      .write_en(par_done_reg1115_write_en),
      .clk(clk),
      .out(par_done_reg1115_out),
      .done(par_done_reg1115_done)
  );
  
  std_reg #(1) par_done_reg1116 (
      .in(par_done_reg1116_in),
      .write_en(par_done_reg1116_write_en),
      .clk(clk),
      .out(par_done_reg1116_out),
      .done(par_done_reg1116_done)
  );
  
  std_reg #(1) par_done_reg1117 (
      .in(par_done_reg1117_in),
      .write_en(par_done_reg1117_write_en),
      .clk(clk),
      .out(par_done_reg1117_out),
      .done(par_done_reg1117_done)
  );
  
  std_reg #(1) par_done_reg1118 (
      .in(par_done_reg1118_in),
      .write_en(par_done_reg1118_write_en),
      .clk(clk),
      .out(par_done_reg1118_out),
      .done(par_done_reg1118_done)
  );
  
  std_reg #(1) par_done_reg1119 (
      .in(par_done_reg1119_in),
      .write_en(par_done_reg1119_write_en),
      .clk(clk),
      .out(par_done_reg1119_out),
      .done(par_done_reg1119_done)
  );
  
  std_reg #(1) par_done_reg1120 (
      .in(par_done_reg1120_in),
      .write_en(par_done_reg1120_write_en),
      .clk(clk),
      .out(par_done_reg1120_out),
      .done(par_done_reg1120_done)
  );
  
  std_reg #(1) par_done_reg1121 (
      .in(par_done_reg1121_in),
      .write_en(par_done_reg1121_write_en),
      .clk(clk),
      .out(par_done_reg1121_out),
      .done(par_done_reg1121_done)
  );
  
  std_reg #(1) par_done_reg1122 (
      .in(par_done_reg1122_in),
      .write_en(par_done_reg1122_write_en),
      .clk(clk),
      .out(par_done_reg1122_out),
      .done(par_done_reg1122_done)
  );
  
  std_reg #(1) par_done_reg1123 (
      .in(par_done_reg1123_in),
      .write_en(par_done_reg1123_write_en),
      .clk(clk),
      .out(par_done_reg1123_out),
      .done(par_done_reg1123_done)
  );
  
  std_reg #(1) par_done_reg1124 (
      .in(par_done_reg1124_in),
      .write_en(par_done_reg1124_write_en),
      .clk(clk),
      .out(par_done_reg1124_out),
      .done(par_done_reg1124_done)
  );
  
  std_reg #(1) par_done_reg1125 (
      .in(par_done_reg1125_in),
      .write_en(par_done_reg1125_write_en),
      .clk(clk),
      .out(par_done_reg1125_out),
      .done(par_done_reg1125_done)
  );
  
  std_reg #(1) par_done_reg1126 (
      .in(par_done_reg1126_in),
      .write_en(par_done_reg1126_write_en),
      .clk(clk),
      .out(par_done_reg1126_out),
      .done(par_done_reg1126_done)
  );
  
  std_reg #(1) par_done_reg1127 (
      .in(par_done_reg1127_in),
      .write_en(par_done_reg1127_write_en),
      .clk(clk),
      .out(par_done_reg1127_out),
      .done(par_done_reg1127_done)
  );
  
  std_reg #(1) par_done_reg1128 (
      .in(par_done_reg1128_in),
      .write_en(par_done_reg1128_write_en),
      .clk(clk),
      .out(par_done_reg1128_out),
      .done(par_done_reg1128_done)
  );
  
  std_reg #(1) par_done_reg1129 (
      .in(par_done_reg1129_in),
      .write_en(par_done_reg1129_write_en),
      .clk(clk),
      .out(par_done_reg1129_out),
      .done(par_done_reg1129_done)
  );
  
  std_reg #(1) par_done_reg1130 (
      .in(par_done_reg1130_in),
      .write_en(par_done_reg1130_write_en),
      .clk(clk),
      .out(par_done_reg1130_out),
      .done(par_done_reg1130_done)
  );
  
  std_reg #(1) par_done_reg1131 (
      .in(par_done_reg1131_in),
      .write_en(par_done_reg1131_write_en),
      .clk(clk),
      .out(par_done_reg1131_out),
      .done(par_done_reg1131_done)
  );
  
  std_reg #(1) par_done_reg1132 (
      .in(par_done_reg1132_in),
      .write_en(par_done_reg1132_write_en),
      .clk(clk),
      .out(par_done_reg1132_out),
      .done(par_done_reg1132_done)
  );
  
  std_reg #(1) par_done_reg1133 (
      .in(par_done_reg1133_in),
      .write_en(par_done_reg1133_write_en),
      .clk(clk),
      .out(par_done_reg1133_out),
      .done(par_done_reg1133_done)
  );
  
  std_reg #(1) par_done_reg1134 (
      .in(par_done_reg1134_in),
      .write_en(par_done_reg1134_write_en),
      .clk(clk),
      .out(par_done_reg1134_out),
      .done(par_done_reg1134_done)
  );
  
  std_reg #(1) par_done_reg1135 (
      .in(par_done_reg1135_in),
      .write_en(par_done_reg1135_write_en),
      .clk(clk),
      .out(par_done_reg1135_out),
      .done(par_done_reg1135_done)
  );
  
  std_reg #(1) par_done_reg1136 (
      .in(par_done_reg1136_in),
      .write_en(par_done_reg1136_write_en),
      .clk(clk),
      .out(par_done_reg1136_out),
      .done(par_done_reg1136_done)
  );
  
  std_reg #(1) par_done_reg1137 (
      .in(par_done_reg1137_in),
      .write_en(par_done_reg1137_write_en),
      .clk(clk),
      .out(par_done_reg1137_out),
      .done(par_done_reg1137_done)
  );
  
  std_reg #(1) par_done_reg1138 (
      .in(par_done_reg1138_in),
      .write_en(par_done_reg1138_write_en),
      .clk(clk),
      .out(par_done_reg1138_out),
      .done(par_done_reg1138_done)
  );
  
  std_reg #(1) par_done_reg1139 (
      .in(par_done_reg1139_in),
      .write_en(par_done_reg1139_write_en),
      .clk(clk),
      .out(par_done_reg1139_out),
      .done(par_done_reg1139_done)
  );
  
  std_reg #(1) par_done_reg1140 (
      .in(par_done_reg1140_in),
      .write_en(par_done_reg1140_write_en),
      .clk(clk),
      .out(par_done_reg1140_out),
      .done(par_done_reg1140_done)
  );
  
  std_reg #(1) par_done_reg1141 (
      .in(par_done_reg1141_in),
      .write_en(par_done_reg1141_write_en),
      .clk(clk),
      .out(par_done_reg1141_out),
      .done(par_done_reg1141_done)
  );
  
  std_reg #(1) par_reset27 (
      .in(par_reset27_in),
      .write_en(par_reset27_write_en),
      .clk(clk),
      .out(par_reset27_out),
      .done(par_reset27_done)
  );
  
  std_reg #(1) par_done_reg1142 (
      .in(par_done_reg1142_in),
      .write_en(par_done_reg1142_write_en),
      .clk(clk),
      .out(par_done_reg1142_out),
      .done(par_done_reg1142_done)
  );
  
  std_reg #(1) par_done_reg1143 (
      .in(par_done_reg1143_in),
      .write_en(par_done_reg1143_write_en),
      .clk(clk),
      .out(par_done_reg1143_out),
      .done(par_done_reg1143_done)
  );
  
  std_reg #(1) par_done_reg1144 (
      .in(par_done_reg1144_in),
      .write_en(par_done_reg1144_write_en),
      .clk(clk),
      .out(par_done_reg1144_out),
      .done(par_done_reg1144_done)
  );
  
  std_reg #(1) par_done_reg1145 (
      .in(par_done_reg1145_in),
      .write_en(par_done_reg1145_write_en),
      .clk(clk),
      .out(par_done_reg1145_out),
      .done(par_done_reg1145_done)
  );
  
  std_reg #(1) par_done_reg1146 (
      .in(par_done_reg1146_in),
      .write_en(par_done_reg1146_write_en),
      .clk(clk),
      .out(par_done_reg1146_out),
      .done(par_done_reg1146_done)
  );
  
  std_reg #(1) par_done_reg1147 (
      .in(par_done_reg1147_in),
      .write_en(par_done_reg1147_write_en),
      .clk(clk),
      .out(par_done_reg1147_out),
      .done(par_done_reg1147_done)
  );
  
  std_reg #(1) par_done_reg1148 (
      .in(par_done_reg1148_in),
      .write_en(par_done_reg1148_write_en),
      .clk(clk),
      .out(par_done_reg1148_out),
      .done(par_done_reg1148_done)
  );
  
  std_reg #(1) par_done_reg1149 (
      .in(par_done_reg1149_in),
      .write_en(par_done_reg1149_write_en),
      .clk(clk),
      .out(par_done_reg1149_out),
      .done(par_done_reg1149_done)
  );
  
  std_reg #(1) par_done_reg1150 (
      .in(par_done_reg1150_in),
      .write_en(par_done_reg1150_write_en),
      .clk(clk),
      .out(par_done_reg1150_out),
      .done(par_done_reg1150_done)
  );
  
  std_reg #(1) par_done_reg1151 (
      .in(par_done_reg1151_in),
      .write_en(par_done_reg1151_write_en),
      .clk(clk),
      .out(par_done_reg1151_out),
      .done(par_done_reg1151_done)
  );
  
  std_reg #(1) par_done_reg1152 (
      .in(par_done_reg1152_in),
      .write_en(par_done_reg1152_write_en),
      .clk(clk),
      .out(par_done_reg1152_out),
      .done(par_done_reg1152_done)
  );
  
  std_reg #(1) par_done_reg1153 (
      .in(par_done_reg1153_in),
      .write_en(par_done_reg1153_write_en),
      .clk(clk),
      .out(par_done_reg1153_out),
      .done(par_done_reg1153_done)
  );
  
  std_reg #(1) par_done_reg1154 (
      .in(par_done_reg1154_in),
      .write_en(par_done_reg1154_write_en),
      .clk(clk),
      .out(par_done_reg1154_out),
      .done(par_done_reg1154_done)
  );
  
  std_reg #(1) par_done_reg1155 (
      .in(par_done_reg1155_in),
      .write_en(par_done_reg1155_write_en),
      .clk(clk),
      .out(par_done_reg1155_out),
      .done(par_done_reg1155_done)
  );
  
  std_reg #(1) par_done_reg1156 (
      .in(par_done_reg1156_in),
      .write_en(par_done_reg1156_write_en),
      .clk(clk),
      .out(par_done_reg1156_out),
      .done(par_done_reg1156_done)
  );
  
  std_reg #(1) par_done_reg1157 (
      .in(par_done_reg1157_in),
      .write_en(par_done_reg1157_write_en),
      .clk(clk),
      .out(par_done_reg1157_out),
      .done(par_done_reg1157_done)
  );
  
  std_reg #(1) par_done_reg1158 (
      .in(par_done_reg1158_in),
      .write_en(par_done_reg1158_write_en),
      .clk(clk),
      .out(par_done_reg1158_out),
      .done(par_done_reg1158_done)
  );
  
  std_reg #(1) par_done_reg1159 (
      .in(par_done_reg1159_in),
      .write_en(par_done_reg1159_write_en),
      .clk(clk),
      .out(par_done_reg1159_out),
      .done(par_done_reg1159_done)
  );
  
  std_reg #(1) par_done_reg1160 (
      .in(par_done_reg1160_in),
      .write_en(par_done_reg1160_write_en),
      .clk(clk),
      .out(par_done_reg1160_out),
      .done(par_done_reg1160_done)
  );
  
  std_reg #(1) par_done_reg1161 (
      .in(par_done_reg1161_in),
      .write_en(par_done_reg1161_write_en),
      .clk(clk),
      .out(par_done_reg1161_out),
      .done(par_done_reg1161_done)
  );
  
  std_reg #(1) par_done_reg1162 (
      .in(par_done_reg1162_in),
      .write_en(par_done_reg1162_write_en),
      .clk(clk),
      .out(par_done_reg1162_out),
      .done(par_done_reg1162_done)
  );
  
  std_reg #(1) par_done_reg1163 (
      .in(par_done_reg1163_in),
      .write_en(par_done_reg1163_write_en),
      .clk(clk),
      .out(par_done_reg1163_out),
      .done(par_done_reg1163_done)
  );
  
  std_reg #(1) par_done_reg1164 (
      .in(par_done_reg1164_in),
      .write_en(par_done_reg1164_write_en),
      .clk(clk),
      .out(par_done_reg1164_out),
      .done(par_done_reg1164_done)
  );
  
  std_reg #(1) par_done_reg1165 (
      .in(par_done_reg1165_in),
      .write_en(par_done_reg1165_write_en),
      .clk(clk),
      .out(par_done_reg1165_out),
      .done(par_done_reg1165_done)
  );
  
  std_reg #(1) par_done_reg1166 (
      .in(par_done_reg1166_in),
      .write_en(par_done_reg1166_write_en),
      .clk(clk),
      .out(par_done_reg1166_out),
      .done(par_done_reg1166_done)
  );
  
  std_reg #(1) par_done_reg1167 (
      .in(par_done_reg1167_in),
      .write_en(par_done_reg1167_write_en),
      .clk(clk),
      .out(par_done_reg1167_out),
      .done(par_done_reg1167_done)
  );
  
  std_reg #(1) par_done_reg1168 (
      .in(par_done_reg1168_in),
      .write_en(par_done_reg1168_write_en),
      .clk(clk),
      .out(par_done_reg1168_out),
      .done(par_done_reg1168_done)
  );
  
  std_reg #(1) par_done_reg1169 (
      .in(par_done_reg1169_in),
      .write_en(par_done_reg1169_write_en),
      .clk(clk),
      .out(par_done_reg1169_out),
      .done(par_done_reg1169_done)
  );
  
  std_reg #(1) par_done_reg1170 (
      .in(par_done_reg1170_in),
      .write_en(par_done_reg1170_write_en),
      .clk(clk),
      .out(par_done_reg1170_out),
      .done(par_done_reg1170_done)
  );
  
  std_reg #(1) par_done_reg1171 (
      .in(par_done_reg1171_in),
      .write_en(par_done_reg1171_write_en),
      .clk(clk),
      .out(par_done_reg1171_out),
      .done(par_done_reg1171_done)
  );
  
  std_reg #(1) par_done_reg1172 (
      .in(par_done_reg1172_in),
      .write_en(par_done_reg1172_write_en),
      .clk(clk),
      .out(par_done_reg1172_out),
      .done(par_done_reg1172_done)
  );
  
  std_reg #(1) par_done_reg1173 (
      .in(par_done_reg1173_in),
      .write_en(par_done_reg1173_write_en),
      .clk(clk),
      .out(par_done_reg1173_out),
      .done(par_done_reg1173_done)
  );
  
  std_reg #(1) par_done_reg1174 (
      .in(par_done_reg1174_in),
      .write_en(par_done_reg1174_write_en),
      .clk(clk),
      .out(par_done_reg1174_out),
      .done(par_done_reg1174_done)
  );
  
  std_reg #(1) par_done_reg1175 (
      .in(par_done_reg1175_in),
      .write_en(par_done_reg1175_write_en),
      .clk(clk),
      .out(par_done_reg1175_out),
      .done(par_done_reg1175_done)
  );
  
  std_reg #(1) par_done_reg1176 (
      .in(par_done_reg1176_in),
      .write_en(par_done_reg1176_write_en),
      .clk(clk),
      .out(par_done_reg1176_out),
      .done(par_done_reg1176_done)
  );
  
  std_reg #(1) par_done_reg1177 (
      .in(par_done_reg1177_in),
      .write_en(par_done_reg1177_write_en),
      .clk(clk),
      .out(par_done_reg1177_out),
      .done(par_done_reg1177_done)
  );
  
  std_reg #(1) par_done_reg1178 (
      .in(par_done_reg1178_in),
      .write_en(par_done_reg1178_write_en),
      .clk(clk),
      .out(par_done_reg1178_out),
      .done(par_done_reg1178_done)
  );
  
  std_reg #(1) par_done_reg1179 (
      .in(par_done_reg1179_in),
      .write_en(par_done_reg1179_write_en),
      .clk(clk),
      .out(par_done_reg1179_out),
      .done(par_done_reg1179_done)
  );
  
  std_reg #(1) par_done_reg1180 (
      .in(par_done_reg1180_in),
      .write_en(par_done_reg1180_write_en),
      .clk(clk),
      .out(par_done_reg1180_out),
      .done(par_done_reg1180_done)
  );
  
  std_reg #(1) par_done_reg1181 (
      .in(par_done_reg1181_in),
      .write_en(par_done_reg1181_write_en),
      .clk(clk),
      .out(par_done_reg1181_out),
      .done(par_done_reg1181_done)
  );
  
  std_reg #(1) par_done_reg1182 (
      .in(par_done_reg1182_in),
      .write_en(par_done_reg1182_write_en),
      .clk(clk),
      .out(par_done_reg1182_out),
      .done(par_done_reg1182_done)
  );
  
  std_reg #(1) par_done_reg1183 (
      .in(par_done_reg1183_in),
      .write_en(par_done_reg1183_write_en),
      .clk(clk),
      .out(par_done_reg1183_out),
      .done(par_done_reg1183_done)
  );
  
  std_reg #(1) par_done_reg1184 (
      .in(par_done_reg1184_in),
      .write_en(par_done_reg1184_write_en),
      .clk(clk),
      .out(par_done_reg1184_out),
      .done(par_done_reg1184_done)
  );
  
  std_reg #(1) par_done_reg1185 (
      .in(par_done_reg1185_in),
      .write_en(par_done_reg1185_write_en),
      .clk(clk),
      .out(par_done_reg1185_out),
      .done(par_done_reg1185_done)
  );
  
  std_reg #(1) par_done_reg1186 (
      .in(par_done_reg1186_in),
      .write_en(par_done_reg1186_write_en),
      .clk(clk),
      .out(par_done_reg1186_out),
      .done(par_done_reg1186_done)
  );
  
  std_reg #(1) par_done_reg1187 (
      .in(par_done_reg1187_in),
      .write_en(par_done_reg1187_write_en),
      .clk(clk),
      .out(par_done_reg1187_out),
      .done(par_done_reg1187_done)
  );
  
  std_reg #(1) par_done_reg1188 (
      .in(par_done_reg1188_in),
      .write_en(par_done_reg1188_write_en),
      .clk(clk),
      .out(par_done_reg1188_out),
      .done(par_done_reg1188_done)
  );
  
  std_reg #(1) par_done_reg1189 (
      .in(par_done_reg1189_in),
      .write_en(par_done_reg1189_write_en),
      .clk(clk),
      .out(par_done_reg1189_out),
      .done(par_done_reg1189_done)
  );
  
  std_reg #(1) par_done_reg1190 (
      .in(par_done_reg1190_in),
      .write_en(par_done_reg1190_write_en),
      .clk(clk),
      .out(par_done_reg1190_out),
      .done(par_done_reg1190_done)
  );
  
  std_reg #(1) par_done_reg1191 (
      .in(par_done_reg1191_in),
      .write_en(par_done_reg1191_write_en),
      .clk(clk),
      .out(par_done_reg1191_out),
      .done(par_done_reg1191_done)
  );
  
  std_reg #(1) par_reset28 (
      .in(par_reset28_in),
      .write_en(par_reset28_write_en),
      .clk(clk),
      .out(par_reset28_out),
      .done(par_reset28_done)
  );
  
  std_reg #(1) par_done_reg1192 (
      .in(par_done_reg1192_in),
      .write_en(par_done_reg1192_write_en),
      .clk(clk),
      .out(par_done_reg1192_out),
      .done(par_done_reg1192_done)
  );
  
  std_reg #(1) par_done_reg1193 (
      .in(par_done_reg1193_in),
      .write_en(par_done_reg1193_write_en),
      .clk(clk),
      .out(par_done_reg1193_out),
      .done(par_done_reg1193_done)
  );
  
  std_reg #(1) par_done_reg1194 (
      .in(par_done_reg1194_in),
      .write_en(par_done_reg1194_write_en),
      .clk(clk),
      .out(par_done_reg1194_out),
      .done(par_done_reg1194_done)
  );
  
  std_reg #(1) par_done_reg1195 (
      .in(par_done_reg1195_in),
      .write_en(par_done_reg1195_write_en),
      .clk(clk),
      .out(par_done_reg1195_out),
      .done(par_done_reg1195_done)
  );
  
  std_reg #(1) par_done_reg1196 (
      .in(par_done_reg1196_in),
      .write_en(par_done_reg1196_write_en),
      .clk(clk),
      .out(par_done_reg1196_out),
      .done(par_done_reg1196_done)
  );
  
  std_reg #(1) par_done_reg1197 (
      .in(par_done_reg1197_in),
      .write_en(par_done_reg1197_write_en),
      .clk(clk),
      .out(par_done_reg1197_out),
      .done(par_done_reg1197_done)
  );
  
  std_reg #(1) par_done_reg1198 (
      .in(par_done_reg1198_in),
      .write_en(par_done_reg1198_write_en),
      .clk(clk),
      .out(par_done_reg1198_out),
      .done(par_done_reg1198_done)
  );
  
  std_reg #(1) par_done_reg1199 (
      .in(par_done_reg1199_in),
      .write_en(par_done_reg1199_write_en),
      .clk(clk),
      .out(par_done_reg1199_out),
      .done(par_done_reg1199_done)
  );
  
  std_reg #(1) par_done_reg1200 (
      .in(par_done_reg1200_in),
      .write_en(par_done_reg1200_write_en),
      .clk(clk),
      .out(par_done_reg1200_out),
      .done(par_done_reg1200_done)
  );
  
  std_reg #(1) par_done_reg1201 (
      .in(par_done_reg1201_in),
      .write_en(par_done_reg1201_write_en),
      .clk(clk),
      .out(par_done_reg1201_out),
      .done(par_done_reg1201_done)
  );
  
  std_reg #(1) par_done_reg1202 (
      .in(par_done_reg1202_in),
      .write_en(par_done_reg1202_write_en),
      .clk(clk),
      .out(par_done_reg1202_out),
      .done(par_done_reg1202_done)
  );
  
  std_reg #(1) par_done_reg1203 (
      .in(par_done_reg1203_in),
      .write_en(par_done_reg1203_write_en),
      .clk(clk),
      .out(par_done_reg1203_out),
      .done(par_done_reg1203_done)
  );
  
  std_reg #(1) par_done_reg1204 (
      .in(par_done_reg1204_in),
      .write_en(par_done_reg1204_write_en),
      .clk(clk),
      .out(par_done_reg1204_out),
      .done(par_done_reg1204_done)
  );
  
  std_reg #(1) par_done_reg1205 (
      .in(par_done_reg1205_in),
      .write_en(par_done_reg1205_write_en),
      .clk(clk),
      .out(par_done_reg1205_out),
      .done(par_done_reg1205_done)
  );
  
  std_reg #(1) par_done_reg1206 (
      .in(par_done_reg1206_in),
      .write_en(par_done_reg1206_write_en),
      .clk(clk),
      .out(par_done_reg1206_out),
      .done(par_done_reg1206_done)
  );
  
  std_reg #(1) par_done_reg1207 (
      .in(par_done_reg1207_in),
      .write_en(par_done_reg1207_write_en),
      .clk(clk),
      .out(par_done_reg1207_out),
      .done(par_done_reg1207_done)
  );
  
  std_reg #(1) par_done_reg1208 (
      .in(par_done_reg1208_in),
      .write_en(par_done_reg1208_write_en),
      .clk(clk),
      .out(par_done_reg1208_out),
      .done(par_done_reg1208_done)
  );
  
  std_reg #(1) par_done_reg1209 (
      .in(par_done_reg1209_in),
      .write_en(par_done_reg1209_write_en),
      .clk(clk),
      .out(par_done_reg1209_out),
      .done(par_done_reg1209_done)
  );
  
  std_reg #(1) par_done_reg1210 (
      .in(par_done_reg1210_in),
      .write_en(par_done_reg1210_write_en),
      .clk(clk),
      .out(par_done_reg1210_out),
      .done(par_done_reg1210_done)
  );
  
  std_reg #(1) par_done_reg1211 (
      .in(par_done_reg1211_in),
      .write_en(par_done_reg1211_write_en),
      .clk(clk),
      .out(par_done_reg1211_out),
      .done(par_done_reg1211_done)
  );
  
  std_reg #(1) par_done_reg1212 (
      .in(par_done_reg1212_in),
      .write_en(par_done_reg1212_write_en),
      .clk(clk),
      .out(par_done_reg1212_out),
      .done(par_done_reg1212_done)
  );
  
  std_reg #(1) par_done_reg1213 (
      .in(par_done_reg1213_in),
      .write_en(par_done_reg1213_write_en),
      .clk(clk),
      .out(par_done_reg1213_out),
      .done(par_done_reg1213_done)
  );
  
  std_reg #(1) par_done_reg1214 (
      .in(par_done_reg1214_in),
      .write_en(par_done_reg1214_write_en),
      .clk(clk),
      .out(par_done_reg1214_out),
      .done(par_done_reg1214_done)
  );
  
  std_reg #(1) par_done_reg1215 (
      .in(par_done_reg1215_in),
      .write_en(par_done_reg1215_write_en),
      .clk(clk),
      .out(par_done_reg1215_out),
      .done(par_done_reg1215_done)
  );
  
  std_reg #(1) par_done_reg1216 (
      .in(par_done_reg1216_in),
      .write_en(par_done_reg1216_write_en),
      .clk(clk),
      .out(par_done_reg1216_out),
      .done(par_done_reg1216_done)
  );
  
  std_reg #(1) par_done_reg1217 (
      .in(par_done_reg1217_in),
      .write_en(par_done_reg1217_write_en),
      .clk(clk),
      .out(par_done_reg1217_out),
      .done(par_done_reg1217_done)
  );
  
  std_reg #(1) par_done_reg1218 (
      .in(par_done_reg1218_in),
      .write_en(par_done_reg1218_write_en),
      .clk(clk),
      .out(par_done_reg1218_out),
      .done(par_done_reg1218_done)
  );
  
  std_reg #(1) par_done_reg1219 (
      .in(par_done_reg1219_in),
      .write_en(par_done_reg1219_write_en),
      .clk(clk),
      .out(par_done_reg1219_out),
      .done(par_done_reg1219_done)
  );
  
  std_reg #(1) par_done_reg1220 (
      .in(par_done_reg1220_in),
      .write_en(par_done_reg1220_write_en),
      .clk(clk),
      .out(par_done_reg1220_out),
      .done(par_done_reg1220_done)
  );
  
  std_reg #(1) par_done_reg1221 (
      .in(par_done_reg1221_in),
      .write_en(par_done_reg1221_write_en),
      .clk(clk),
      .out(par_done_reg1221_out),
      .done(par_done_reg1221_done)
  );
  
  std_reg #(1) par_done_reg1222 (
      .in(par_done_reg1222_in),
      .write_en(par_done_reg1222_write_en),
      .clk(clk),
      .out(par_done_reg1222_out),
      .done(par_done_reg1222_done)
  );
  
  std_reg #(1) par_done_reg1223 (
      .in(par_done_reg1223_in),
      .write_en(par_done_reg1223_write_en),
      .clk(clk),
      .out(par_done_reg1223_out),
      .done(par_done_reg1223_done)
  );
  
  std_reg #(1) par_done_reg1224 (
      .in(par_done_reg1224_in),
      .write_en(par_done_reg1224_write_en),
      .clk(clk),
      .out(par_done_reg1224_out),
      .done(par_done_reg1224_done)
  );
  
  std_reg #(1) par_done_reg1225 (
      .in(par_done_reg1225_in),
      .write_en(par_done_reg1225_write_en),
      .clk(clk),
      .out(par_done_reg1225_out),
      .done(par_done_reg1225_done)
  );
  
  std_reg #(1) par_done_reg1226 (
      .in(par_done_reg1226_in),
      .write_en(par_done_reg1226_write_en),
      .clk(clk),
      .out(par_done_reg1226_out),
      .done(par_done_reg1226_done)
  );
  
  std_reg #(1) par_done_reg1227 (
      .in(par_done_reg1227_in),
      .write_en(par_done_reg1227_write_en),
      .clk(clk),
      .out(par_done_reg1227_out),
      .done(par_done_reg1227_done)
  );
  
  std_reg #(1) par_done_reg1228 (
      .in(par_done_reg1228_in),
      .write_en(par_done_reg1228_write_en),
      .clk(clk),
      .out(par_done_reg1228_out),
      .done(par_done_reg1228_done)
  );
  
  std_reg #(1) par_done_reg1229 (
      .in(par_done_reg1229_in),
      .write_en(par_done_reg1229_write_en),
      .clk(clk),
      .out(par_done_reg1229_out),
      .done(par_done_reg1229_done)
  );
  
  std_reg #(1) par_done_reg1230 (
      .in(par_done_reg1230_in),
      .write_en(par_done_reg1230_write_en),
      .clk(clk),
      .out(par_done_reg1230_out),
      .done(par_done_reg1230_done)
  );
  
  std_reg #(1) par_done_reg1231 (
      .in(par_done_reg1231_in),
      .write_en(par_done_reg1231_write_en),
      .clk(clk),
      .out(par_done_reg1231_out),
      .done(par_done_reg1231_done)
  );
  
  std_reg #(1) par_done_reg1232 (
      .in(par_done_reg1232_in),
      .write_en(par_done_reg1232_write_en),
      .clk(clk),
      .out(par_done_reg1232_out),
      .done(par_done_reg1232_done)
  );
  
  std_reg #(1) par_done_reg1233 (
      .in(par_done_reg1233_in),
      .write_en(par_done_reg1233_write_en),
      .clk(clk),
      .out(par_done_reg1233_out),
      .done(par_done_reg1233_done)
  );
  
  std_reg #(1) par_done_reg1234 (
      .in(par_done_reg1234_in),
      .write_en(par_done_reg1234_write_en),
      .clk(clk),
      .out(par_done_reg1234_out),
      .done(par_done_reg1234_done)
  );
  
  std_reg #(1) par_done_reg1235 (
      .in(par_done_reg1235_in),
      .write_en(par_done_reg1235_write_en),
      .clk(clk),
      .out(par_done_reg1235_out),
      .done(par_done_reg1235_done)
  );
  
  std_reg #(1) par_done_reg1236 (
      .in(par_done_reg1236_in),
      .write_en(par_done_reg1236_write_en),
      .clk(clk),
      .out(par_done_reg1236_out),
      .done(par_done_reg1236_done)
  );
  
  std_reg #(1) par_done_reg1237 (
      .in(par_done_reg1237_in),
      .write_en(par_done_reg1237_write_en),
      .clk(clk),
      .out(par_done_reg1237_out),
      .done(par_done_reg1237_done)
  );
  
  std_reg #(1) par_done_reg1238 (
      .in(par_done_reg1238_in),
      .write_en(par_done_reg1238_write_en),
      .clk(clk),
      .out(par_done_reg1238_out),
      .done(par_done_reg1238_done)
  );
  
  std_reg #(1) par_done_reg1239 (
      .in(par_done_reg1239_in),
      .write_en(par_done_reg1239_write_en),
      .clk(clk),
      .out(par_done_reg1239_out),
      .done(par_done_reg1239_done)
  );
  
  std_reg #(1) par_done_reg1240 (
      .in(par_done_reg1240_in),
      .write_en(par_done_reg1240_write_en),
      .clk(clk),
      .out(par_done_reg1240_out),
      .done(par_done_reg1240_done)
  );
  
  std_reg #(1) par_done_reg1241 (
      .in(par_done_reg1241_in),
      .write_en(par_done_reg1241_write_en),
      .clk(clk),
      .out(par_done_reg1241_out),
      .done(par_done_reg1241_done)
  );
  
  std_reg #(1) par_done_reg1242 (
      .in(par_done_reg1242_in),
      .write_en(par_done_reg1242_write_en),
      .clk(clk),
      .out(par_done_reg1242_out),
      .done(par_done_reg1242_done)
  );
  
  std_reg #(1) par_done_reg1243 (
      .in(par_done_reg1243_in),
      .write_en(par_done_reg1243_write_en),
      .clk(clk),
      .out(par_done_reg1243_out),
      .done(par_done_reg1243_done)
  );
  
  std_reg #(1) par_done_reg1244 (
      .in(par_done_reg1244_in),
      .write_en(par_done_reg1244_write_en),
      .clk(clk),
      .out(par_done_reg1244_out),
      .done(par_done_reg1244_done)
  );
  
  std_reg #(1) par_done_reg1245 (
      .in(par_done_reg1245_in),
      .write_en(par_done_reg1245_write_en),
      .clk(clk),
      .out(par_done_reg1245_out),
      .done(par_done_reg1245_done)
  );
  
  std_reg #(1) par_done_reg1246 (
      .in(par_done_reg1246_in),
      .write_en(par_done_reg1246_write_en),
      .clk(clk),
      .out(par_done_reg1246_out),
      .done(par_done_reg1246_done)
  );
  
  std_reg #(1) par_done_reg1247 (
      .in(par_done_reg1247_in),
      .write_en(par_done_reg1247_write_en),
      .clk(clk),
      .out(par_done_reg1247_out),
      .done(par_done_reg1247_done)
  );
  
  std_reg #(1) par_done_reg1248 (
      .in(par_done_reg1248_in),
      .write_en(par_done_reg1248_write_en),
      .clk(clk),
      .out(par_done_reg1248_out),
      .done(par_done_reg1248_done)
  );
  
  std_reg #(1) par_done_reg1249 (
      .in(par_done_reg1249_in),
      .write_en(par_done_reg1249_write_en),
      .clk(clk),
      .out(par_done_reg1249_out),
      .done(par_done_reg1249_done)
  );
  
  std_reg #(1) par_done_reg1250 (
      .in(par_done_reg1250_in),
      .write_en(par_done_reg1250_write_en),
      .clk(clk),
      .out(par_done_reg1250_out),
      .done(par_done_reg1250_done)
  );
  
  std_reg #(1) par_done_reg1251 (
      .in(par_done_reg1251_in),
      .write_en(par_done_reg1251_write_en),
      .clk(clk),
      .out(par_done_reg1251_out),
      .done(par_done_reg1251_done)
  );
  
  std_reg #(1) par_done_reg1252 (
      .in(par_done_reg1252_in),
      .write_en(par_done_reg1252_write_en),
      .clk(clk),
      .out(par_done_reg1252_out),
      .done(par_done_reg1252_done)
  );
  
  std_reg #(1) par_done_reg1253 (
      .in(par_done_reg1253_in),
      .write_en(par_done_reg1253_write_en),
      .clk(clk),
      .out(par_done_reg1253_out),
      .done(par_done_reg1253_done)
  );
  
  std_reg #(1) par_done_reg1254 (
      .in(par_done_reg1254_in),
      .write_en(par_done_reg1254_write_en),
      .clk(clk),
      .out(par_done_reg1254_out),
      .done(par_done_reg1254_done)
  );
  
  std_reg #(1) par_done_reg1255 (
      .in(par_done_reg1255_in),
      .write_en(par_done_reg1255_write_en),
      .clk(clk),
      .out(par_done_reg1255_out),
      .done(par_done_reg1255_done)
  );
  
  std_reg #(1) par_done_reg1256 (
      .in(par_done_reg1256_in),
      .write_en(par_done_reg1256_write_en),
      .clk(clk),
      .out(par_done_reg1256_out),
      .done(par_done_reg1256_done)
  );
  
  std_reg #(1) par_done_reg1257 (
      .in(par_done_reg1257_in),
      .write_en(par_done_reg1257_write_en),
      .clk(clk),
      .out(par_done_reg1257_out),
      .done(par_done_reg1257_done)
  );
  
  std_reg #(1) par_done_reg1258 (
      .in(par_done_reg1258_in),
      .write_en(par_done_reg1258_write_en),
      .clk(clk),
      .out(par_done_reg1258_out),
      .done(par_done_reg1258_done)
  );
  
  std_reg #(1) par_done_reg1259 (
      .in(par_done_reg1259_in),
      .write_en(par_done_reg1259_write_en),
      .clk(clk),
      .out(par_done_reg1259_out),
      .done(par_done_reg1259_done)
  );
  
  std_reg #(1) par_done_reg1260 (
      .in(par_done_reg1260_in),
      .write_en(par_done_reg1260_write_en),
      .clk(clk),
      .out(par_done_reg1260_out),
      .done(par_done_reg1260_done)
  );
  
  std_reg #(1) par_done_reg1261 (
      .in(par_done_reg1261_in),
      .write_en(par_done_reg1261_write_en),
      .clk(clk),
      .out(par_done_reg1261_out),
      .done(par_done_reg1261_done)
  );
  
  std_reg #(1) par_done_reg1262 (
      .in(par_done_reg1262_in),
      .write_en(par_done_reg1262_write_en),
      .clk(clk),
      .out(par_done_reg1262_out),
      .done(par_done_reg1262_done)
  );
  
  std_reg #(1) par_done_reg1263 (
      .in(par_done_reg1263_in),
      .write_en(par_done_reg1263_write_en),
      .clk(clk),
      .out(par_done_reg1263_out),
      .done(par_done_reg1263_done)
  );
  
  std_reg #(1) par_done_reg1264 (
      .in(par_done_reg1264_in),
      .write_en(par_done_reg1264_write_en),
      .clk(clk),
      .out(par_done_reg1264_out),
      .done(par_done_reg1264_done)
  );
  
  std_reg #(1) par_done_reg1265 (
      .in(par_done_reg1265_in),
      .write_en(par_done_reg1265_write_en),
      .clk(clk),
      .out(par_done_reg1265_out),
      .done(par_done_reg1265_done)
  );
  
  std_reg #(1) par_done_reg1266 (
      .in(par_done_reg1266_in),
      .write_en(par_done_reg1266_write_en),
      .clk(clk),
      .out(par_done_reg1266_out),
      .done(par_done_reg1266_done)
  );
  
  std_reg #(1) par_done_reg1267 (
      .in(par_done_reg1267_in),
      .write_en(par_done_reg1267_write_en),
      .clk(clk),
      .out(par_done_reg1267_out),
      .done(par_done_reg1267_done)
  );
  
  std_reg #(1) par_done_reg1268 (
      .in(par_done_reg1268_in),
      .write_en(par_done_reg1268_write_en),
      .clk(clk),
      .out(par_done_reg1268_out),
      .done(par_done_reg1268_done)
  );
  
  std_reg #(1) par_done_reg1269 (
      .in(par_done_reg1269_in),
      .write_en(par_done_reg1269_write_en),
      .clk(clk),
      .out(par_done_reg1269_out),
      .done(par_done_reg1269_done)
  );
  
  std_reg #(1) par_done_reg1270 (
      .in(par_done_reg1270_in),
      .write_en(par_done_reg1270_write_en),
      .clk(clk),
      .out(par_done_reg1270_out),
      .done(par_done_reg1270_done)
  );
  
  std_reg #(1) par_done_reg1271 (
      .in(par_done_reg1271_in),
      .write_en(par_done_reg1271_write_en),
      .clk(clk),
      .out(par_done_reg1271_out),
      .done(par_done_reg1271_done)
  );
  
  std_reg #(1) par_done_reg1272 (
      .in(par_done_reg1272_in),
      .write_en(par_done_reg1272_write_en),
      .clk(clk),
      .out(par_done_reg1272_out),
      .done(par_done_reg1272_done)
  );
  
  std_reg #(1) par_done_reg1273 (
      .in(par_done_reg1273_in),
      .write_en(par_done_reg1273_write_en),
      .clk(clk),
      .out(par_done_reg1273_out),
      .done(par_done_reg1273_done)
  );
  
  std_reg #(1) par_done_reg1274 (
      .in(par_done_reg1274_in),
      .write_en(par_done_reg1274_write_en),
      .clk(clk),
      .out(par_done_reg1274_out),
      .done(par_done_reg1274_done)
  );
  
  std_reg #(1) par_done_reg1275 (
      .in(par_done_reg1275_in),
      .write_en(par_done_reg1275_write_en),
      .clk(clk),
      .out(par_done_reg1275_out),
      .done(par_done_reg1275_done)
  );
  
  std_reg #(1) par_reset29 (
      .in(par_reset29_in),
      .write_en(par_reset29_write_en),
      .clk(clk),
      .out(par_reset29_out),
      .done(par_reset29_done)
  );
  
  std_reg #(1) par_done_reg1276 (
      .in(par_done_reg1276_in),
      .write_en(par_done_reg1276_write_en),
      .clk(clk),
      .out(par_done_reg1276_out),
      .done(par_done_reg1276_done)
  );
  
  std_reg #(1) par_done_reg1277 (
      .in(par_done_reg1277_in),
      .write_en(par_done_reg1277_write_en),
      .clk(clk),
      .out(par_done_reg1277_out),
      .done(par_done_reg1277_done)
  );
  
  std_reg #(1) par_done_reg1278 (
      .in(par_done_reg1278_in),
      .write_en(par_done_reg1278_write_en),
      .clk(clk),
      .out(par_done_reg1278_out),
      .done(par_done_reg1278_done)
  );
  
  std_reg #(1) par_done_reg1279 (
      .in(par_done_reg1279_in),
      .write_en(par_done_reg1279_write_en),
      .clk(clk),
      .out(par_done_reg1279_out),
      .done(par_done_reg1279_done)
  );
  
  std_reg #(1) par_done_reg1280 (
      .in(par_done_reg1280_in),
      .write_en(par_done_reg1280_write_en),
      .clk(clk),
      .out(par_done_reg1280_out),
      .done(par_done_reg1280_done)
  );
  
  std_reg #(1) par_done_reg1281 (
      .in(par_done_reg1281_in),
      .write_en(par_done_reg1281_write_en),
      .clk(clk),
      .out(par_done_reg1281_out),
      .done(par_done_reg1281_done)
  );
  
  std_reg #(1) par_done_reg1282 (
      .in(par_done_reg1282_in),
      .write_en(par_done_reg1282_write_en),
      .clk(clk),
      .out(par_done_reg1282_out),
      .done(par_done_reg1282_done)
  );
  
  std_reg #(1) par_done_reg1283 (
      .in(par_done_reg1283_in),
      .write_en(par_done_reg1283_write_en),
      .clk(clk),
      .out(par_done_reg1283_out),
      .done(par_done_reg1283_done)
  );
  
  std_reg #(1) par_done_reg1284 (
      .in(par_done_reg1284_in),
      .write_en(par_done_reg1284_write_en),
      .clk(clk),
      .out(par_done_reg1284_out),
      .done(par_done_reg1284_done)
  );
  
  std_reg #(1) par_done_reg1285 (
      .in(par_done_reg1285_in),
      .write_en(par_done_reg1285_write_en),
      .clk(clk),
      .out(par_done_reg1285_out),
      .done(par_done_reg1285_done)
  );
  
  std_reg #(1) par_done_reg1286 (
      .in(par_done_reg1286_in),
      .write_en(par_done_reg1286_write_en),
      .clk(clk),
      .out(par_done_reg1286_out),
      .done(par_done_reg1286_done)
  );
  
  std_reg #(1) par_done_reg1287 (
      .in(par_done_reg1287_in),
      .write_en(par_done_reg1287_write_en),
      .clk(clk),
      .out(par_done_reg1287_out),
      .done(par_done_reg1287_done)
  );
  
  std_reg #(1) par_done_reg1288 (
      .in(par_done_reg1288_in),
      .write_en(par_done_reg1288_write_en),
      .clk(clk),
      .out(par_done_reg1288_out),
      .done(par_done_reg1288_done)
  );
  
  std_reg #(1) par_done_reg1289 (
      .in(par_done_reg1289_in),
      .write_en(par_done_reg1289_write_en),
      .clk(clk),
      .out(par_done_reg1289_out),
      .done(par_done_reg1289_done)
  );
  
  std_reg #(1) par_done_reg1290 (
      .in(par_done_reg1290_in),
      .write_en(par_done_reg1290_write_en),
      .clk(clk),
      .out(par_done_reg1290_out),
      .done(par_done_reg1290_done)
  );
  
  std_reg #(1) par_done_reg1291 (
      .in(par_done_reg1291_in),
      .write_en(par_done_reg1291_write_en),
      .clk(clk),
      .out(par_done_reg1291_out),
      .done(par_done_reg1291_done)
  );
  
  std_reg #(1) par_done_reg1292 (
      .in(par_done_reg1292_in),
      .write_en(par_done_reg1292_write_en),
      .clk(clk),
      .out(par_done_reg1292_out),
      .done(par_done_reg1292_done)
  );
  
  std_reg #(1) par_done_reg1293 (
      .in(par_done_reg1293_in),
      .write_en(par_done_reg1293_write_en),
      .clk(clk),
      .out(par_done_reg1293_out),
      .done(par_done_reg1293_done)
  );
  
  std_reg #(1) par_done_reg1294 (
      .in(par_done_reg1294_in),
      .write_en(par_done_reg1294_write_en),
      .clk(clk),
      .out(par_done_reg1294_out),
      .done(par_done_reg1294_done)
  );
  
  std_reg #(1) par_done_reg1295 (
      .in(par_done_reg1295_in),
      .write_en(par_done_reg1295_write_en),
      .clk(clk),
      .out(par_done_reg1295_out),
      .done(par_done_reg1295_done)
  );
  
  std_reg #(1) par_done_reg1296 (
      .in(par_done_reg1296_in),
      .write_en(par_done_reg1296_write_en),
      .clk(clk),
      .out(par_done_reg1296_out),
      .done(par_done_reg1296_done)
  );
  
  std_reg #(1) par_done_reg1297 (
      .in(par_done_reg1297_in),
      .write_en(par_done_reg1297_write_en),
      .clk(clk),
      .out(par_done_reg1297_out),
      .done(par_done_reg1297_done)
  );
  
  std_reg #(1) par_done_reg1298 (
      .in(par_done_reg1298_in),
      .write_en(par_done_reg1298_write_en),
      .clk(clk),
      .out(par_done_reg1298_out),
      .done(par_done_reg1298_done)
  );
  
  std_reg #(1) par_done_reg1299 (
      .in(par_done_reg1299_in),
      .write_en(par_done_reg1299_write_en),
      .clk(clk),
      .out(par_done_reg1299_out),
      .done(par_done_reg1299_done)
  );
  
  std_reg #(1) par_done_reg1300 (
      .in(par_done_reg1300_in),
      .write_en(par_done_reg1300_write_en),
      .clk(clk),
      .out(par_done_reg1300_out),
      .done(par_done_reg1300_done)
  );
  
  std_reg #(1) par_done_reg1301 (
      .in(par_done_reg1301_in),
      .write_en(par_done_reg1301_write_en),
      .clk(clk),
      .out(par_done_reg1301_out),
      .done(par_done_reg1301_done)
  );
  
  std_reg #(1) par_done_reg1302 (
      .in(par_done_reg1302_in),
      .write_en(par_done_reg1302_write_en),
      .clk(clk),
      .out(par_done_reg1302_out),
      .done(par_done_reg1302_done)
  );
  
  std_reg #(1) par_done_reg1303 (
      .in(par_done_reg1303_in),
      .write_en(par_done_reg1303_write_en),
      .clk(clk),
      .out(par_done_reg1303_out),
      .done(par_done_reg1303_done)
  );
  
  std_reg #(1) par_done_reg1304 (
      .in(par_done_reg1304_in),
      .write_en(par_done_reg1304_write_en),
      .clk(clk),
      .out(par_done_reg1304_out),
      .done(par_done_reg1304_done)
  );
  
  std_reg #(1) par_done_reg1305 (
      .in(par_done_reg1305_in),
      .write_en(par_done_reg1305_write_en),
      .clk(clk),
      .out(par_done_reg1305_out),
      .done(par_done_reg1305_done)
  );
  
  std_reg #(1) par_done_reg1306 (
      .in(par_done_reg1306_in),
      .write_en(par_done_reg1306_write_en),
      .clk(clk),
      .out(par_done_reg1306_out),
      .done(par_done_reg1306_done)
  );
  
  std_reg #(1) par_done_reg1307 (
      .in(par_done_reg1307_in),
      .write_en(par_done_reg1307_write_en),
      .clk(clk),
      .out(par_done_reg1307_out),
      .done(par_done_reg1307_done)
  );
  
  std_reg #(1) par_done_reg1308 (
      .in(par_done_reg1308_in),
      .write_en(par_done_reg1308_write_en),
      .clk(clk),
      .out(par_done_reg1308_out),
      .done(par_done_reg1308_done)
  );
  
  std_reg #(1) par_done_reg1309 (
      .in(par_done_reg1309_in),
      .write_en(par_done_reg1309_write_en),
      .clk(clk),
      .out(par_done_reg1309_out),
      .done(par_done_reg1309_done)
  );
  
  std_reg #(1) par_done_reg1310 (
      .in(par_done_reg1310_in),
      .write_en(par_done_reg1310_write_en),
      .clk(clk),
      .out(par_done_reg1310_out),
      .done(par_done_reg1310_done)
  );
  
  std_reg #(1) par_done_reg1311 (
      .in(par_done_reg1311_in),
      .write_en(par_done_reg1311_write_en),
      .clk(clk),
      .out(par_done_reg1311_out),
      .done(par_done_reg1311_done)
  );
  
  std_reg #(1) par_done_reg1312 (
      .in(par_done_reg1312_in),
      .write_en(par_done_reg1312_write_en),
      .clk(clk),
      .out(par_done_reg1312_out),
      .done(par_done_reg1312_done)
  );
  
  std_reg #(1) par_done_reg1313 (
      .in(par_done_reg1313_in),
      .write_en(par_done_reg1313_write_en),
      .clk(clk),
      .out(par_done_reg1313_out),
      .done(par_done_reg1313_done)
  );
  
  std_reg #(1) par_done_reg1314 (
      .in(par_done_reg1314_in),
      .write_en(par_done_reg1314_write_en),
      .clk(clk),
      .out(par_done_reg1314_out),
      .done(par_done_reg1314_done)
  );
  
  std_reg #(1) par_done_reg1315 (
      .in(par_done_reg1315_in),
      .write_en(par_done_reg1315_write_en),
      .clk(clk),
      .out(par_done_reg1315_out),
      .done(par_done_reg1315_done)
  );
  
  std_reg #(1) par_done_reg1316 (
      .in(par_done_reg1316_in),
      .write_en(par_done_reg1316_write_en),
      .clk(clk),
      .out(par_done_reg1316_out),
      .done(par_done_reg1316_done)
  );
  
  std_reg #(1) par_done_reg1317 (
      .in(par_done_reg1317_in),
      .write_en(par_done_reg1317_write_en),
      .clk(clk),
      .out(par_done_reg1317_out),
      .done(par_done_reg1317_done)
  );
  
  std_reg #(1) par_done_reg1318 (
      .in(par_done_reg1318_in),
      .write_en(par_done_reg1318_write_en),
      .clk(clk),
      .out(par_done_reg1318_out),
      .done(par_done_reg1318_done)
  );
  
  std_reg #(1) par_done_reg1319 (
      .in(par_done_reg1319_in),
      .write_en(par_done_reg1319_write_en),
      .clk(clk),
      .out(par_done_reg1319_out),
      .done(par_done_reg1319_done)
  );
  
  std_reg #(1) par_reset30 (
      .in(par_reset30_in),
      .write_en(par_reset30_write_en),
      .clk(clk),
      .out(par_reset30_out),
      .done(par_reset30_done)
  );
  
  std_reg #(1) par_done_reg1320 (
      .in(par_done_reg1320_in),
      .write_en(par_done_reg1320_write_en),
      .clk(clk),
      .out(par_done_reg1320_out),
      .done(par_done_reg1320_done)
  );
  
  std_reg #(1) par_done_reg1321 (
      .in(par_done_reg1321_in),
      .write_en(par_done_reg1321_write_en),
      .clk(clk),
      .out(par_done_reg1321_out),
      .done(par_done_reg1321_done)
  );
  
  std_reg #(1) par_done_reg1322 (
      .in(par_done_reg1322_in),
      .write_en(par_done_reg1322_write_en),
      .clk(clk),
      .out(par_done_reg1322_out),
      .done(par_done_reg1322_done)
  );
  
  std_reg #(1) par_done_reg1323 (
      .in(par_done_reg1323_in),
      .write_en(par_done_reg1323_write_en),
      .clk(clk),
      .out(par_done_reg1323_out),
      .done(par_done_reg1323_done)
  );
  
  std_reg #(1) par_done_reg1324 (
      .in(par_done_reg1324_in),
      .write_en(par_done_reg1324_write_en),
      .clk(clk),
      .out(par_done_reg1324_out),
      .done(par_done_reg1324_done)
  );
  
  std_reg #(1) par_done_reg1325 (
      .in(par_done_reg1325_in),
      .write_en(par_done_reg1325_write_en),
      .clk(clk),
      .out(par_done_reg1325_out),
      .done(par_done_reg1325_done)
  );
  
  std_reg #(1) par_done_reg1326 (
      .in(par_done_reg1326_in),
      .write_en(par_done_reg1326_write_en),
      .clk(clk),
      .out(par_done_reg1326_out),
      .done(par_done_reg1326_done)
  );
  
  std_reg #(1) par_done_reg1327 (
      .in(par_done_reg1327_in),
      .write_en(par_done_reg1327_write_en),
      .clk(clk),
      .out(par_done_reg1327_out),
      .done(par_done_reg1327_done)
  );
  
  std_reg #(1) par_done_reg1328 (
      .in(par_done_reg1328_in),
      .write_en(par_done_reg1328_write_en),
      .clk(clk),
      .out(par_done_reg1328_out),
      .done(par_done_reg1328_done)
  );
  
  std_reg #(1) par_done_reg1329 (
      .in(par_done_reg1329_in),
      .write_en(par_done_reg1329_write_en),
      .clk(clk),
      .out(par_done_reg1329_out),
      .done(par_done_reg1329_done)
  );
  
  std_reg #(1) par_done_reg1330 (
      .in(par_done_reg1330_in),
      .write_en(par_done_reg1330_write_en),
      .clk(clk),
      .out(par_done_reg1330_out),
      .done(par_done_reg1330_done)
  );
  
  std_reg #(1) par_done_reg1331 (
      .in(par_done_reg1331_in),
      .write_en(par_done_reg1331_write_en),
      .clk(clk),
      .out(par_done_reg1331_out),
      .done(par_done_reg1331_done)
  );
  
  std_reg #(1) par_done_reg1332 (
      .in(par_done_reg1332_in),
      .write_en(par_done_reg1332_write_en),
      .clk(clk),
      .out(par_done_reg1332_out),
      .done(par_done_reg1332_done)
  );
  
  std_reg #(1) par_done_reg1333 (
      .in(par_done_reg1333_in),
      .write_en(par_done_reg1333_write_en),
      .clk(clk),
      .out(par_done_reg1333_out),
      .done(par_done_reg1333_done)
  );
  
  std_reg #(1) par_done_reg1334 (
      .in(par_done_reg1334_in),
      .write_en(par_done_reg1334_write_en),
      .clk(clk),
      .out(par_done_reg1334_out),
      .done(par_done_reg1334_done)
  );
  
  std_reg #(1) par_done_reg1335 (
      .in(par_done_reg1335_in),
      .write_en(par_done_reg1335_write_en),
      .clk(clk),
      .out(par_done_reg1335_out),
      .done(par_done_reg1335_done)
  );
  
  std_reg #(1) par_done_reg1336 (
      .in(par_done_reg1336_in),
      .write_en(par_done_reg1336_write_en),
      .clk(clk),
      .out(par_done_reg1336_out),
      .done(par_done_reg1336_done)
  );
  
  std_reg #(1) par_done_reg1337 (
      .in(par_done_reg1337_in),
      .write_en(par_done_reg1337_write_en),
      .clk(clk),
      .out(par_done_reg1337_out),
      .done(par_done_reg1337_done)
  );
  
  std_reg #(1) par_done_reg1338 (
      .in(par_done_reg1338_in),
      .write_en(par_done_reg1338_write_en),
      .clk(clk),
      .out(par_done_reg1338_out),
      .done(par_done_reg1338_done)
  );
  
  std_reg #(1) par_done_reg1339 (
      .in(par_done_reg1339_in),
      .write_en(par_done_reg1339_write_en),
      .clk(clk),
      .out(par_done_reg1339_out),
      .done(par_done_reg1339_done)
  );
  
  std_reg #(1) par_done_reg1340 (
      .in(par_done_reg1340_in),
      .write_en(par_done_reg1340_write_en),
      .clk(clk),
      .out(par_done_reg1340_out),
      .done(par_done_reg1340_done)
  );
  
  std_reg #(1) par_done_reg1341 (
      .in(par_done_reg1341_in),
      .write_en(par_done_reg1341_write_en),
      .clk(clk),
      .out(par_done_reg1341_out),
      .done(par_done_reg1341_done)
  );
  
  std_reg #(1) par_done_reg1342 (
      .in(par_done_reg1342_in),
      .write_en(par_done_reg1342_write_en),
      .clk(clk),
      .out(par_done_reg1342_out),
      .done(par_done_reg1342_done)
  );
  
  std_reg #(1) par_done_reg1343 (
      .in(par_done_reg1343_in),
      .write_en(par_done_reg1343_write_en),
      .clk(clk),
      .out(par_done_reg1343_out),
      .done(par_done_reg1343_done)
  );
  
  std_reg #(1) par_done_reg1344 (
      .in(par_done_reg1344_in),
      .write_en(par_done_reg1344_write_en),
      .clk(clk),
      .out(par_done_reg1344_out),
      .done(par_done_reg1344_done)
  );
  
  std_reg #(1) par_done_reg1345 (
      .in(par_done_reg1345_in),
      .write_en(par_done_reg1345_write_en),
      .clk(clk),
      .out(par_done_reg1345_out),
      .done(par_done_reg1345_done)
  );
  
  std_reg #(1) par_done_reg1346 (
      .in(par_done_reg1346_in),
      .write_en(par_done_reg1346_write_en),
      .clk(clk),
      .out(par_done_reg1346_out),
      .done(par_done_reg1346_done)
  );
  
  std_reg #(1) par_done_reg1347 (
      .in(par_done_reg1347_in),
      .write_en(par_done_reg1347_write_en),
      .clk(clk),
      .out(par_done_reg1347_out),
      .done(par_done_reg1347_done)
  );
  
  std_reg #(1) par_done_reg1348 (
      .in(par_done_reg1348_in),
      .write_en(par_done_reg1348_write_en),
      .clk(clk),
      .out(par_done_reg1348_out),
      .done(par_done_reg1348_done)
  );
  
  std_reg #(1) par_done_reg1349 (
      .in(par_done_reg1349_in),
      .write_en(par_done_reg1349_write_en),
      .clk(clk),
      .out(par_done_reg1349_out),
      .done(par_done_reg1349_done)
  );
  
  std_reg #(1) par_done_reg1350 (
      .in(par_done_reg1350_in),
      .write_en(par_done_reg1350_write_en),
      .clk(clk),
      .out(par_done_reg1350_out),
      .done(par_done_reg1350_done)
  );
  
  std_reg #(1) par_done_reg1351 (
      .in(par_done_reg1351_in),
      .write_en(par_done_reg1351_write_en),
      .clk(clk),
      .out(par_done_reg1351_out),
      .done(par_done_reg1351_done)
  );
  
  std_reg #(1) par_done_reg1352 (
      .in(par_done_reg1352_in),
      .write_en(par_done_reg1352_write_en),
      .clk(clk),
      .out(par_done_reg1352_out),
      .done(par_done_reg1352_done)
  );
  
  std_reg #(1) par_done_reg1353 (
      .in(par_done_reg1353_in),
      .write_en(par_done_reg1353_write_en),
      .clk(clk),
      .out(par_done_reg1353_out),
      .done(par_done_reg1353_done)
  );
  
  std_reg #(1) par_done_reg1354 (
      .in(par_done_reg1354_in),
      .write_en(par_done_reg1354_write_en),
      .clk(clk),
      .out(par_done_reg1354_out),
      .done(par_done_reg1354_done)
  );
  
  std_reg #(1) par_done_reg1355 (
      .in(par_done_reg1355_in),
      .write_en(par_done_reg1355_write_en),
      .clk(clk),
      .out(par_done_reg1355_out),
      .done(par_done_reg1355_done)
  );
  
  std_reg #(1) par_done_reg1356 (
      .in(par_done_reg1356_in),
      .write_en(par_done_reg1356_write_en),
      .clk(clk),
      .out(par_done_reg1356_out),
      .done(par_done_reg1356_done)
  );
  
  std_reg #(1) par_done_reg1357 (
      .in(par_done_reg1357_in),
      .write_en(par_done_reg1357_write_en),
      .clk(clk),
      .out(par_done_reg1357_out),
      .done(par_done_reg1357_done)
  );
  
  std_reg #(1) par_done_reg1358 (
      .in(par_done_reg1358_in),
      .write_en(par_done_reg1358_write_en),
      .clk(clk),
      .out(par_done_reg1358_out),
      .done(par_done_reg1358_done)
  );
  
  std_reg #(1) par_done_reg1359 (
      .in(par_done_reg1359_in),
      .write_en(par_done_reg1359_write_en),
      .clk(clk),
      .out(par_done_reg1359_out),
      .done(par_done_reg1359_done)
  );
  
  std_reg #(1) par_done_reg1360 (
      .in(par_done_reg1360_in),
      .write_en(par_done_reg1360_write_en),
      .clk(clk),
      .out(par_done_reg1360_out),
      .done(par_done_reg1360_done)
  );
  
  std_reg #(1) par_done_reg1361 (
      .in(par_done_reg1361_in),
      .write_en(par_done_reg1361_write_en),
      .clk(clk),
      .out(par_done_reg1361_out),
      .done(par_done_reg1361_done)
  );
  
  std_reg #(1) par_done_reg1362 (
      .in(par_done_reg1362_in),
      .write_en(par_done_reg1362_write_en),
      .clk(clk),
      .out(par_done_reg1362_out),
      .done(par_done_reg1362_done)
  );
  
  std_reg #(1) par_done_reg1363 (
      .in(par_done_reg1363_in),
      .write_en(par_done_reg1363_write_en),
      .clk(clk),
      .out(par_done_reg1363_out),
      .done(par_done_reg1363_done)
  );
  
  std_reg #(1) par_done_reg1364 (
      .in(par_done_reg1364_in),
      .write_en(par_done_reg1364_write_en),
      .clk(clk),
      .out(par_done_reg1364_out),
      .done(par_done_reg1364_done)
  );
  
  std_reg #(1) par_done_reg1365 (
      .in(par_done_reg1365_in),
      .write_en(par_done_reg1365_write_en),
      .clk(clk),
      .out(par_done_reg1365_out),
      .done(par_done_reg1365_done)
  );
  
  std_reg #(1) par_done_reg1366 (
      .in(par_done_reg1366_in),
      .write_en(par_done_reg1366_write_en),
      .clk(clk),
      .out(par_done_reg1366_out),
      .done(par_done_reg1366_done)
  );
  
  std_reg #(1) par_done_reg1367 (
      .in(par_done_reg1367_in),
      .write_en(par_done_reg1367_write_en),
      .clk(clk),
      .out(par_done_reg1367_out),
      .done(par_done_reg1367_done)
  );
  
  std_reg #(1) par_done_reg1368 (
      .in(par_done_reg1368_in),
      .write_en(par_done_reg1368_write_en),
      .clk(clk),
      .out(par_done_reg1368_out),
      .done(par_done_reg1368_done)
  );
  
  std_reg #(1) par_done_reg1369 (
      .in(par_done_reg1369_in),
      .write_en(par_done_reg1369_write_en),
      .clk(clk),
      .out(par_done_reg1369_out),
      .done(par_done_reg1369_done)
  );
  
  std_reg #(1) par_done_reg1370 (
      .in(par_done_reg1370_in),
      .write_en(par_done_reg1370_write_en),
      .clk(clk),
      .out(par_done_reg1370_out),
      .done(par_done_reg1370_done)
  );
  
  std_reg #(1) par_done_reg1371 (
      .in(par_done_reg1371_in),
      .write_en(par_done_reg1371_write_en),
      .clk(clk),
      .out(par_done_reg1371_out),
      .done(par_done_reg1371_done)
  );
  
  std_reg #(1) par_done_reg1372 (
      .in(par_done_reg1372_in),
      .write_en(par_done_reg1372_write_en),
      .clk(clk),
      .out(par_done_reg1372_out),
      .done(par_done_reg1372_done)
  );
  
  std_reg #(1) par_done_reg1373 (
      .in(par_done_reg1373_in),
      .write_en(par_done_reg1373_write_en),
      .clk(clk),
      .out(par_done_reg1373_out),
      .done(par_done_reg1373_done)
  );
  
  std_reg #(1) par_done_reg1374 (
      .in(par_done_reg1374_in),
      .write_en(par_done_reg1374_write_en),
      .clk(clk),
      .out(par_done_reg1374_out),
      .done(par_done_reg1374_done)
  );
  
  std_reg #(1) par_done_reg1375 (
      .in(par_done_reg1375_in),
      .write_en(par_done_reg1375_write_en),
      .clk(clk),
      .out(par_done_reg1375_out),
      .done(par_done_reg1375_done)
  );
  
  std_reg #(1) par_done_reg1376 (
      .in(par_done_reg1376_in),
      .write_en(par_done_reg1376_write_en),
      .clk(clk),
      .out(par_done_reg1376_out),
      .done(par_done_reg1376_done)
  );
  
  std_reg #(1) par_done_reg1377 (
      .in(par_done_reg1377_in),
      .write_en(par_done_reg1377_write_en),
      .clk(clk),
      .out(par_done_reg1377_out),
      .done(par_done_reg1377_done)
  );
  
  std_reg #(1) par_done_reg1378 (
      .in(par_done_reg1378_in),
      .write_en(par_done_reg1378_write_en),
      .clk(clk),
      .out(par_done_reg1378_out),
      .done(par_done_reg1378_done)
  );
  
  std_reg #(1) par_done_reg1379 (
      .in(par_done_reg1379_in),
      .write_en(par_done_reg1379_write_en),
      .clk(clk),
      .out(par_done_reg1379_out),
      .done(par_done_reg1379_done)
  );
  
  std_reg #(1) par_done_reg1380 (
      .in(par_done_reg1380_in),
      .write_en(par_done_reg1380_write_en),
      .clk(clk),
      .out(par_done_reg1380_out),
      .done(par_done_reg1380_done)
  );
  
  std_reg #(1) par_done_reg1381 (
      .in(par_done_reg1381_in),
      .write_en(par_done_reg1381_write_en),
      .clk(clk),
      .out(par_done_reg1381_out),
      .done(par_done_reg1381_done)
  );
  
  std_reg #(1) par_done_reg1382 (
      .in(par_done_reg1382_in),
      .write_en(par_done_reg1382_write_en),
      .clk(clk),
      .out(par_done_reg1382_out),
      .done(par_done_reg1382_done)
  );
  
  std_reg #(1) par_done_reg1383 (
      .in(par_done_reg1383_in),
      .write_en(par_done_reg1383_write_en),
      .clk(clk),
      .out(par_done_reg1383_out),
      .done(par_done_reg1383_done)
  );
  
  std_reg #(1) par_done_reg1384 (
      .in(par_done_reg1384_in),
      .write_en(par_done_reg1384_write_en),
      .clk(clk),
      .out(par_done_reg1384_out),
      .done(par_done_reg1384_done)
  );
  
  std_reg #(1) par_done_reg1385 (
      .in(par_done_reg1385_in),
      .write_en(par_done_reg1385_write_en),
      .clk(clk),
      .out(par_done_reg1385_out),
      .done(par_done_reg1385_done)
  );
  
  std_reg #(1) par_done_reg1386 (
      .in(par_done_reg1386_in),
      .write_en(par_done_reg1386_write_en),
      .clk(clk),
      .out(par_done_reg1386_out),
      .done(par_done_reg1386_done)
  );
  
  std_reg #(1) par_done_reg1387 (
      .in(par_done_reg1387_in),
      .write_en(par_done_reg1387_write_en),
      .clk(clk),
      .out(par_done_reg1387_out),
      .done(par_done_reg1387_done)
  );
  
  std_reg #(1) par_done_reg1388 (
      .in(par_done_reg1388_in),
      .write_en(par_done_reg1388_write_en),
      .clk(clk),
      .out(par_done_reg1388_out),
      .done(par_done_reg1388_done)
  );
  
  std_reg #(1) par_done_reg1389 (
      .in(par_done_reg1389_in),
      .write_en(par_done_reg1389_write_en),
      .clk(clk),
      .out(par_done_reg1389_out),
      .done(par_done_reg1389_done)
  );
  
  std_reg #(1) par_done_reg1390 (
      .in(par_done_reg1390_in),
      .write_en(par_done_reg1390_write_en),
      .clk(clk),
      .out(par_done_reg1390_out),
      .done(par_done_reg1390_done)
  );
  
  std_reg #(1) par_done_reg1391 (
      .in(par_done_reg1391_in),
      .write_en(par_done_reg1391_write_en),
      .clk(clk),
      .out(par_done_reg1391_out),
      .done(par_done_reg1391_done)
  );
  
  std_reg #(1) par_reset31 (
      .in(par_reset31_in),
      .write_en(par_reset31_write_en),
      .clk(clk),
      .out(par_reset31_out),
      .done(par_reset31_done)
  );
  
  std_reg #(1) par_done_reg1392 (
      .in(par_done_reg1392_in),
      .write_en(par_done_reg1392_write_en),
      .clk(clk),
      .out(par_done_reg1392_out),
      .done(par_done_reg1392_done)
  );
  
  std_reg #(1) par_done_reg1393 (
      .in(par_done_reg1393_in),
      .write_en(par_done_reg1393_write_en),
      .clk(clk),
      .out(par_done_reg1393_out),
      .done(par_done_reg1393_done)
  );
  
  std_reg #(1) par_done_reg1394 (
      .in(par_done_reg1394_in),
      .write_en(par_done_reg1394_write_en),
      .clk(clk),
      .out(par_done_reg1394_out),
      .done(par_done_reg1394_done)
  );
  
  std_reg #(1) par_done_reg1395 (
      .in(par_done_reg1395_in),
      .write_en(par_done_reg1395_write_en),
      .clk(clk),
      .out(par_done_reg1395_out),
      .done(par_done_reg1395_done)
  );
  
  std_reg #(1) par_done_reg1396 (
      .in(par_done_reg1396_in),
      .write_en(par_done_reg1396_write_en),
      .clk(clk),
      .out(par_done_reg1396_out),
      .done(par_done_reg1396_done)
  );
  
  std_reg #(1) par_done_reg1397 (
      .in(par_done_reg1397_in),
      .write_en(par_done_reg1397_write_en),
      .clk(clk),
      .out(par_done_reg1397_out),
      .done(par_done_reg1397_done)
  );
  
  std_reg #(1) par_done_reg1398 (
      .in(par_done_reg1398_in),
      .write_en(par_done_reg1398_write_en),
      .clk(clk),
      .out(par_done_reg1398_out),
      .done(par_done_reg1398_done)
  );
  
  std_reg #(1) par_done_reg1399 (
      .in(par_done_reg1399_in),
      .write_en(par_done_reg1399_write_en),
      .clk(clk),
      .out(par_done_reg1399_out),
      .done(par_done_reg1399_done)
  );
  
  std_reg #(1) par_done_reg1400 (
      .in(par_done_reg1400_in),
      .write_en(par_done_reg1400_write_en),
      .clk(clk),
      .out(par_done_reg1400_out),
      .done(par_done_reg1400_done)
  );
  
  std_reg #(1) par_done_reg1401 (
      .in(par_done_reg1401_in),
      .write_en(par_done_reg1401_write_en),
      .clk(clk),
      .out(par_done_reg1401_out),
      .done(par_done_reg1401_done)
  );
  
  std_reg #(1) par_done_reg1402 (
      .in(par_done_reg1402_in),
      .write_en(par_done_reg1402_write_en),
      .clk(clk),
      .out(par_done_reg1402_out),
      .done(par_done_reg1402_done)
  );
  
  std_reg #(1) par_done_reg1403 (
      .in(par_done_reg1403_in),
      .write_en(par_done_reg1403_write_en),
      .clk(clk),
      .out(par_done_reg1403_out),
      .done(par_done_reg1403_done)
  );
  
  std_reg #(1) par_done_reg1404 (
      .in(par_done_reg1404_in),
      .write_en(par_done_reg1404_write_en),
      .clk(clk),
      .out(par_done_reg1404_out),
      .done(par_done_reg1404_done)
  );
  
  std_reg #(1) par_done_reg1405 (
      .in(par_done_reg1405_in),
      .write_en(par_done_reg1405_write_en),
      .clk(clk),
      .out(par_done_reg1405_out),
      .done(par_done_reg1405_done)
  );
  
  std_reg #(1) par_done_reg1406 (
      .in(par_done_reg1406_in),
      .write_en(par_done_reg1406_write_en),
      .clk(clk),
      .out(par_done_reg1406_out),
      .done(par_done_reg1406_done)
  );
  
  std_reg #(1) par_done_reg1407 (
      .in(par_done_reg1407_in),
      .write_en(par_done_reg1407_write_en),
      .clk(clk),
      .out(par_done_reg1407_out),
      .done(par_done_reg1407_done)
  );
  
  std_reg #(1) par_done_reg1408 (
      .in(par_done_reg1408_in),
      .write_en(par_done_reg1408_write_en),
      .clk(clk),
      .out(par_done_reg1408_out),
      .done(par_done_reg1408_done)
  );
  
  std_reg #(1) par_done_reg1409 (
      .in(par_done_reg1409_in),
      .write_en(par_done_reg1409_write_en),
      .clk(clk),
      .out(par_done_reg1409_out),
      .done(par_done_reg1409_done)
  );
  
  std_reg #(1) par_done_reg1410 (
      .in(par_done_reg1410_in),
      .write_en(par_done_reg1410_write_en),
      .clk(clk),
      .out(par_done_reg1410_out),
      .done(par_done_reg1410_done)
  );
  
  std_reg #(1) par_done_reg1411 (
      .in(par_done_reg1411_in),
      .write_en(par_done_reg1411_write_en),
      .clk(clk),
      .out(par_done_reg1411_out),
      .done(par_done_reg1411_done)
  );
  
  std_reg #(1) par_done_reg1412 (
      .in(par_done_reg1412_in),
      .write_en(par_done_reg1412_write_en),
      .clk(clk),
      .out(par_done_reg1412_out),
      .done(par_done_reg1412_done)
  );
  
  std_reg #(1) par_done_reg1413 (
      .in(par_done_reg1413_in),
      .write_en(par_done_reg1413_write_en),
      .clk(clk),
      .out(par_done_reg1413_out),
      .done(par_done_reg1413_done)
  );
  
  std_reg #(1) par_done_reg1414 (
      .in(par_done_reg1414_in),
      .write_en(par_done_reg1414_write_en),
      .clk(clk),
      .out(par_done_reg1414_out),
      .done(par_done_reg1414_done)
  );
  
  std_reg #(1) par_done_reg1415 (
      .in(par_done_reg1415_in),
      .write_en(par_done_reg1415_write_en),
      .clk(clk),
      .out(par_done_reg1415_out),
      .done(par_done_reg1415_done)
  );
  
  std_reg #(1) par_done_reg1416 (
      .in(par_done_reg1416_in),
      .write_en(par_done_reg1416_write_en),
      .clk(clk),
      .out(par_done_reg1416_out),
      .done(par_done_reg1416_done)
  );
  
  std_reg #(1) par_done_reg1417 (
      .in(par_done_reg1417_in),
      .write_en(par_done_reg1417_write_en),
      .clk(clk),
      .out(par_done_reg1417_out),
      .done(par_done_reg1417_done)
  );
  
  std_reg #(1) par_done_reg1418 (
      .in(par_done_reg1418_in),
      .write_en(par_done_reg1418_write_en),
      .clk(clk),
      .out(par_done_reg1418_out),
      .done(par_done_reg1418_done)
  );
  
  std_reg #(1) par_done_reg1419 (
      .in(par_done_reg1419_in),
      .write_en(par_done_reg1419_write_en),
      .clk(clk),
      .out(par_done_reg1419_out),
      .done(par_done_reg1419_done)
  );
  
  std_reg #(1) par_done_reg1420 (
      .in(par_done_reg1420_in),
      .write_en(par_done_reg1420_write_en),
      .clk(clk),
      .out(par_done_reg1420_out),
      .done(par_done_reg1420_done)
  );
  
  std_reg #(1) par_done_reg1421 (
      .in(par_done_reg1421_in),
      .write_en(par_done_reg1421_write_en),
      .clk(clk),
      .out(par_done_reg1421_out),
      .done(par_done_reg1421_done)
  );
  
  std_reg #(1) par_done_reg1422 (
      .in(par_done_reg1422_in),
      .write_en(par_done_reg1422_write_en),
      .clk(clk),
      .out(par_done_reg1422_out),
      .done(par_done_reg1422_done)
  );
  
  std_reg #(1) par_done_reg1423 (
      .in(par_done_reg1423_in),
      .write_en(par_done_reg1423_write_en),
      .clk(clk),
      .out(par_done_reg1423_out),
      .done(par_done_reg1423_done)
  );
  
  std_reg #(1) par_done_reg1424 (
      .in(par_done_reg1424_in),
      .write_en(par_done_reg1424_write_en),
      .clk(clk),
      .out(par_done_reg1424_out),
      .done(par_done_reg1424_done)
  );
  
  std_reg #(1) par_done_reg1425 (
      .in(par_done_reg1425_in),
      .write_en(par_done_reg1425_write_en),
      .clk(clk),
      .out(par_done_reg1425_out),
      .done(par_done_reg1425_done)
  );
  
  std_reg #(1) par_done_reg1426 (
      .in(par_done_reg1426_in),
      .write_en(par_done_reg1426_write_en),
      .clk(clk),
      .out(par_done_reg1426_out),
      .done(par_done_reg1426_done)
  );
  
  std_reg #(1) par_done_reg1427 (
      .in(par_done_reg1427_in),
      .write_en(par_done_reg1427_write_en),
      .clk(clk),
      .out(par_done_reg1427_out),
      .done(par_done_reg1427_done)
  );
  
  std_reg #(1) par_reset32 (
      .in(par_reset32_in),
      .write_en(par_reset32_write_en),
      .clk(clk),
      .out(par_reset32_out),
      .done(par_reset32_done)
  );
  
  std_reg #(1) par_done_reg1428 (
      .in(par_done_reg1428_in),
      .write_en(par_done_reg1428_write_en),
      .clk(clk),
      .out(par_done_reg1428_out),
      .done(par_done_reg1428_done)
  );
  
  std_reg #(1) par_done_reg1429 (
      .in(par_done_reg1429_in),
      .write_en(par_done_reg1429_write_en),
      .clk(clk),
      .out(par_done_reg1429_out),
      .done(par_done_reg1429_done)
  );
  
  std_reg #(1) par_done_reg1430 (
      .in(par_done_reg1430_in),
      .write_en(par_done_reg1430_write_en),
      .clk(clk),
      .out(par_done_reg1430_out),
      .done(par_done_reg1430_done)
  );
  
  std_reg #(1) par_done_reg1431 (
      .in(par_done_reg1431_in),
      .write_en(par_done_reg1431_write_en),
      .clk(clk),
      .out(par_done_reg1431_out),
      .done(par_done_reg1431_done)
  );
  
  std_reg #(1) par_done_reg1432 (
      .in(par_done_reg1432_in),
      .write_en(par_done_reg1432_write_en),
      .clk(clk),
      .out(par_done_reg1432_out),
      .done(par_done_reg1432_done)
  );
  
  std_reg #(1) par_done_reg1433 (
      .in(par_done_reg1433_in),
      .write_en(par_done_reg1433_write_en),
      .clk(clk),
      .out(par_done_reg1433_out),
      .done(par_done_reg1433_done)
  );
  
  std_reg #(1) par_done_reg1434 (
      .in(par_done_reg1434_in),
      .write_en(par_done_reg1434_write_en),
      .clk(clk),
      .out(par_done_reg1434_out),
      .done(par_done_reg1434_done)
  );
  
  std_reg #(1) par_done_reg1435 (
      .in(par_done_reg1435_in),
      .write_en(par_done_reg1435_write_en),
      .clk(clk),
      .out(par_done_reg1435_out),
      .done(par_done_reg1435_done)
  );
  
  std_reg #(1) par_done_reg1436 (
      .in(par_done_reg1436_in),
      .write_en(par_done_reg1436_write_en),
      .clk(clk),
      .out(par_done_reg1436_out),
      .done(par_done_reg1436_done)
  );
  
  std_reg #(1) par_done_reg1437 (
      .in(par_done_reg1437_in),
      .write_en(par_done_reg1437_write_en),
      .clk(clk),
      .out(par_done_reg1437_out),
      .done(par_done_reg1437_done)
  );
  
  std_reg #(1) par_done_reg1438 (
      .in(par_done_reg1438_in),
      .write_en(par_done_reg1438_write_en),
      .clk(clk),
      .out(par_done_reg1438_out),
      .done(par_done_reg1438_done)
  );
  
  std_reg #(1) par_done_reg1439 (
      .in(par_done_reg1439_in),
      .write_en(par_done_reg1439_write_en),
      .clk(clk),
      .out(par_done_reg1439_out),
      .done(par_done_reg1439_done)
  );
  
  std_reg #(1) par_done_reg1440 (
      .in(par_done_reg1440_in),
      .write_en(par_done_reg1440_write_en),
      .clk(clk),
      .out(par_done_reg1440_out),
      .done(par_done_reg1440_done)
  );
  
  std_reg #(1) par_done_reg1441 (
      .in(par_done_reg1441_in),
      .write_en(par_done_reg1441_write_en),
      .clk(clk),
      .out(par_done_reg1441_out),
      .done(par_done_reg1441_done)
  );
  
  std_reg #(1) par_done_reg1442 (
      .in(par_done_reg1442_in),
      .write_en(par_done_reg1442_write_en),
      .clk(clk),
      .out(par_done_reg1442_out),
      .done(par_done_reg1442_done)
  );
  
  std_reg #(1) par_done_reg1443 (
      .in(par_done_reg1443_in),
      .write_en(par_done_reg1443_write_en),
      .clk(clk),
      .out(par_done_reg1443_out),
      .done(par_done_reg1443_done)
  );
  
  std_reg #(1) par_done_reg1444 (
      .in(par_done_reg1444_in),
      .write_en(par_done_reg1444_write_en),
      .clk(clk),
      .out(par_done_reg1444_out),
      .done(par_done_reg1444_done)
  );
  
  std_reg #(1) par_done_reg1445 (
      .in(par_done_reg1445_in),
      .write_en(par_done_reg1445_write_en),
      .clk(clk),
      .out(par_done_reg1445_out),
      .done(par_done_reg1445_done)
  );
  
  std_reg #(1) par_done_reg1446 (
      .in(par_done_reg1446_in),
      .write_en(par_done_reg1446_write_en),
      .clk(clk),
      .out(par_done_reg1446_out),
      .done(par_done_reg1446_done)
  );
  
  std_reg #(1) par_done_reg1447 (
      .in(par_done_reg1447_in),
      .write_en(par_done_reg1447_write_en),
      .clk(clk),
      .out(par_done_reg1447_out),
      .done(par_done_reg1447_done)
  );
  
  std_reg #(1) par_done_reg1448 (
      .in(par_done_reg1448_in),
      .write_en(par_done_reg1448_write_en),
      .clk(clk),
      .out(par_done_reg1448_out),
      .done(par_done_reg1448_done)
  );
  
  std_reg #(1) par_done_reg1449 (
      .in(par_done_reg1449_in),
      .write_en(par_done_reg1449_write_en),
      .clk(clk),
      .out(par_done_reg1449_out),
      .done(par_done_reg1449_done)
  );
  
  std_reg #(1) par_done_reg1450 (
      .in(par_done_reg1450_in),
      .write_en(par_done_reg1450_write_en),
      .clk(clk),
      .out(par_done_reg1450_out),
      .done(par_done_reg1450_done)
  );
  
  std_reg #(1) par_done_reg1451 (
      .in(par_done_reg1451_in),
      .write_en(par_done_reg1451_write_en),
      .clk(clk),
      .out(par_done_reg1451_out),
      .done(par_done_reg1451_done)
  );
  
  std_reg #(1) par_done_reg1452 (
      .in(par_done_reg1452_in),
      .write_en(par_done_reg1452_write_en),
      .clk(clk),
      .out(par_done_reg1452_out),
      .done(par_done_reg1452_done)
  );
  
  std_reg #(1) par_done_reg1453 (
      .in(par_done_reg1453_in),
      .write_en(par_done_reg1453_write_en),
      .clk(clk),
      .out(par_done_reg1453_out),
      .done(par_done_reg1453_done)
  );
  
  std_reg #(1) par_done_reg1454 (
      .in(par_done_reg1454_in),
      .write_en(par_done_reg1454_write_en),
      .clk(clk),
      .out(par_done_reg1454_out),
      .done(par_done_reg1454_done)
  );
  
  std_reg #(1) par_done_reg1455 (
      .in(par_done_reg1455_in),
      .write_en(par_done_reg1455_write_en),
      .clk(clk),
      .out(par_done_reg1455_out),
      .done(par_done_reg1455_done)
  );
  
  std_reg #(1) par_done_reg1456 (
      .in(par_done_reg1456_in),
      .write_en(par_done_reg1456_write_en),
      .clk(clk),
      .out(par_done_reg1456_out),
      .done(par_done_reg1456_done)
  );
  
  std_reg #(1) par_done_reg1457 (
      .in(par_done_reg1457_in),
      .write_en(par_done_reg1457_write_en),
      .clk(clk),
      .out(par_done_reg1457_out),
      .done(par_done_reg1457_done)
  );
  
  std_reg #(1) par_done_reg1458 (
      .in(par_done_reg1458_in),
      .write_en(par_done_reg1458_write_en),
      .clk(clk),
      .out(par_done_reg1458_out),
      .done(par_done_reg1458_done)
  );
  
  std_reg #(1) par_done_reg1459 (
      .in(par_done_reg1459_in),
      .write_en(par_done_reg1459_write_en),
      .clk(clk),
      .out(par_done_reg1459_out),
      .done(par_done_reg1459_done)
  );
  
  std_reg #(1) par_done_reg1460 (
      .in(par_done_reg1460_in),
      .write_en(par_done_reg1460_write_en),
      .clk(clk),
      .out(par_done_reg1460_out),
      .done(par_done_reg1460_done)
  );
  
  std_reg #(1) par_done_reg1461 (
      .in(par_done_reg1461_in),
      .write_en(par_done_reg1461_write_en),
      .clk(clk),
      .out(par_done_reg1461_out),
      .done(par_done_reg1461_done)
  );
  
  std_reg #(1) par_done_reg1462 (
      .in(par_done_reg1462_in),
      .write_en(par_done_reg1462_write_en),
      .clk(clk),
      .out(par_done_reg1462_out),
      .done(par_done_reg1462_done)
  );
  
  std_reg #(1) par_done_reg1463 (
      .in(par_done_reg1463_in),
      .write_en(par_done_reg1463_write_en),
      .clk(clk),
      .out(par_done_reg1463_out),
      .done(par_done_reg1463_done)
  );
  
  std_reg #(1) par_done_reg1464 (
      .in(par_done_reg1464_in),
      .write_en(par_done_reg1464_write_en),
      .clk(clk),
      .out(par_done_reg1464_out),
      .done(par_done_reg1464_done)
  );
  
  std_reg #(1) par_done_reg1465 (
      .in(par_done_reg1465_in),
      .write_en(par_done_reg1465_write_en),
      .clk(clk),
      .out(par_done_reg1465_out),
      .done(par_done_reg1465_done)
  );
  
  std_reg #(1) par_done_reg1466 (
      .in(par_done_reg1466_in),
      .write_en(par_done_reg1466_write_en),
      .clk(clk),
      .out(par_done_reg1466_out),
      .done(par_done_reg1466_done)
  );
  
  std_reg #(1) par_done_reg1467 (
      .in(par_done_reg1467_in),
      .write_en(par_done_reg1467_write_en),
      .clk(clk),
      .out(par_done_reg1467_out),
      .done(par_done_reg1467_done)
  );
  
  std_reg #(1) par_done_reg1468 (
      .in(par_done_reg1468_in),
      .write_en(par_done_reg1468_write_en),
      .clk(clk),
      .out(par_done_reg1468_out),
      .done(par_done_reg1468_done)
  );
  
  std_reg #(1) par_done_reg1469 (
      .in(par_done_reg1469_in),
      .write_en(par_done_reg1469_write_en),
      .clk(clk),
      .out(par_done_reg1469_out),
      .done(par_done_reg1469_done)
  );
  
  std_reg #(1) par_done_reg1470 (
      .in(par_done_reg1470_in),
      .write_en(par_done_reg1470_write_en),
      .clk(clk),
      .out(par_done_reg1470_out),
      .done(par_done_reg1470_done)
  );
  
  std_reg #(1) par_done_reg1471 (
      .in(par_done_reg1471_in),
      .write_en(par_done_reg1471_write_en),
      .clk(clk),
      .out(par_done_reg1471_out),
      .done(par_done_reg1471_done)
  );
  
  std_reg #(1) par_done_reg1472 (
      .in(par_done_reg1472_in),
      .write_en(par_done_reg1472_write_en),
      .clk(clk),
      .out(par_done_reg1472_out),
      .done(par_done_reg1472_done)
  );
  
  std_reg #(1) par_done_reg1473 (
      .in(par_done_reg1473_in),
      .write_en(par_done_reg1473_write_en),
      .clk(clk),
      .out(par_done_reg1473_out),
      .done(par_done_reg1473_done)
  );
  
  std_reg #(1) par_done_reg1474 (
      .in(par_done_reg1474_in),
      .write_en(par_done_reg1474_write_en),
      .clk(clk),
      .out(par_done_reg1474_out),
      .done(par_done_reg1474_done)
  );
  
  std_reg #(1) par_done_reg1475 (
      .in(par_done_reg1475_in),
      .write_en(par_done_reg1475_write_en),
      .clk(clk),
      .out(par_done_reg1475_out),
      .done(par_done_reg1475_done)
  );
  
  std_reg #(1) par_done_reg1476 (
      .in(par_done_reg1476_in),
      .write_en(par_done_reg1476_write_en),
      .clk(clk),
      .out(par_done_reg1476_out),
      .done(par_done_reg1476_done)
  );
  
  std_reg #(1) par_done_reg1477 (
      .in(par_done_reg1477_in),
      .write_en(par_done_reg1477_write_en),
      .clk(clk),
      .out(par_done_reg1477_out),
      .done(par_done_reg1477_done)
  );
  
  std_reg #(1) par_done_reg1478 (
      .in(par_done_reg1478_in),
      .write_en(par_done_reg1478_write_en),
      .clk(clk),
      .out(par_done_reg1478_out),
      .done(par_done_reg1478_done)
  );
  
  std_reg #(1) par_done_reg1479 (
      .in(par_done_reg1479_in),
      .write_en(par_done_reg1479_write_en),
      .clk(clk),
      .out(par_done_reg1479_out),
      .done(par_done_reg1479_done)
  );
  
  std_reg #(1) par_done_reg1480 (
      .in(par_done_reg1480_in),
      .write_en(par_done_reg1480_write_en),
      .clk(clk),
      .out(par_done_reg1480_out),
      .done(par_done_reg1480_done)
  );
  
  std_reg #(1) par_done_reg1481 (
      .in(par_done_reg1481_in),
      .write_en(par_done_reg1481_write_en),
      .clk(clk),
      .out(par_done_reg1481_out),
      .done(par_done_reg1481_done)
  );
  
  std_reg #(1) par_done_reg1482 (
      .in(par_done_reg1482_in),
      .write_en(par_done_reg1482_write_en),
      .clk(clk),
      .out(par_done_reg1482_out),
      .done(par_done_reg1482_done)
  );
  
  std_reg #(1) par_done_reg1483 (
      .in(par_done_reg1483_in),
      .write_en(par_done_reg1483_write_en),
      .clk(clk),
      .out(par_done_reg1483_out),
      .done(par_done_reg1483_done)
  );
  
  std_reg #(1) par_reset33 (
      .in(par_reset33_in),
      .write_en(par_reset33_write_en),
      .clk(clk),
      .out(par_reset33_out),
      .done(par_reset33_done)
  );
  
  std_reg #(1) par_done_reg1484 (
      .in(par_done_reg1484_in),
      .write_en(par_done_reg1484_write_en),
      .clk(clk),
      .out(par_done_reg1484_out),
      .done(par_done_reg1484_done)
  );
  
  std_reg #(1) par_done_reg1485 (
      .in(par_done_reg1485_in),
      .write_en(par_done_reg1485_write_en),
      .clk(clk),
      .out(par_done_reg1485_out),
      .done(par_done_reg1485_done)
  );
  
  std_reg #(1) par_done_reg1486 (
      .in(par_done_reg1486_in),
      .write_en(par_done_reg1486_write_en),
      .clk(clk),
      .out(par_done_reg1486_out),
      .done(par_done_reg1486_done)
  );
  
  std_reg #(1) par_done_reg1487 (
      .in(par_done_reg1487_in),
      .write_en(par_done_reg1487_write_en),
      .clk(clk),
      .out(par_done_reg1487_out),
      .done(par_done_reg1487_done)
  );
  
  std_reg #(1) par_done_reg1488 (
      .in(par_done_reg1488_in),
      .write_en(par_done_reg1488_write_en),
      .clk(clk),
      .out(par_done_reg1488_out),
      .done(par_done_reg1488_done)
  );
  
  std_reg #(1) par_done_reg1489 (
      .in(par_done_reg1489_in),
      .write_en(par_done_reg1489_write_en),
      .clk(clk),
      .out(par_done_reg1489_out),
      .done(par_done_reg1489_done)
  );
  
  std_reg #(1) par_done_reg1490 (
      .in(par_done_reg1490_in),
      .write_en(par_done_reg1490_write_en),
      .clk(clk),
      .out(par_done_reg1490_out),
      .done(par_done_reg1490_done)
  );
  
  std_reg #(1) par_done_reg1491 (
      .in(par_done_reg1491_in),
      .write_en(par_done_reg1491_write_en),
      .clk(clk),
      .out(par_done_reg1491_out),
      .done(par_done_reg1491_done)
  );
  
  std_reg #(1) par_done_reg1492 (
      .in(par_done_reg1492_in),
      .write_en(par_done_reg1492_write_en),
      .clk(clk),
      .out(par_done_reg1492_out),
      .done(par_done_reg1492_done)
  );
  
  std_reg #(1) par_done_reg1493 (
      .in(par_done_reg1493_in),
      .write_en(par_done_reg1493_write_en),
      .clk(clk),
      .out(par_done_reg1493_out),
      .done(par_done_reg1493_done)
  );
  
  std_reg #(1) par_done_reg1494 (
      .in(par_done_reg1494_in),
      .write_en(par_done_reg1494_write_en),
      .clk(clk),
      .out(par_done_reg1494_out),
      .done(par_done_reg1494_done)
  );
  
  std_reg #(1) par_done_reg1495 (
      .in(par_done_reg1495_in),
      .write_en(par_done_reg1495_write_en),
      .clk(clk),
      .out(par_done_reg1495_out),
      .done(par_done_reg1495_done)
  );
  
  std_reg #(1) par_done_reg1496 (
      .in(par_done_reg1496_in),
      .write_en(par_done_reg1496_write_en),
      .clk(clk),
      .out(par_done_reg1496_out),
      .done(par_done_reg1496_done)
  );
  
  std_reg #(1) par_done_reg1497 (
      .in(par_done_reg1497_in),
      .write_en(par_done_reg1497_write_en),
      .clk(clk),
      .out(par_done_reg1497_out),
      .done(par_done_reg1497_done)
  );
  
  std_reg #(1) par_done_reg1498 (
      .in(par_done_reg1498_in),
      .write_en(par_done_reg1498_write_en),
      .clk(clk),
      .out(par_done_reg1498_out),
      .done(par_done_reg1498_done)
  );
  
  std_reg #(1) par_done_reg1499 (
      .in(par_done_reg1499_in),
      .write_en(par_done_reg1499_write_en),
      .clk(clk),
      .out(par_done_reg1499_out),
      .done(par_done_reg1499_done)
  );
  
  std_reg #(1) par_done_reg1500 (
      .in(par_done_reg1500_in),
      .write_en(par_done_reg1500_write_en),
      .clk(clk),
      .out(par_done_reg1500_out),
      .done(par_done_reg1500_done)
  );
  
  std_reg #(1) par_done_reg1501 (
      .in(par_done_reg1501_in),
      .write_en(par_done_reg1501_write_en),
      .clk(clk),
      .out(par_done_reg1501_out),
      .done(par_done_reg1501_done)
  );
  
  std_reg #(1) par_done_reg1502 (
      .in(par_done_reg1502_in),
      .write_en(par_done_reg1502_write_en),
      .clk(clk),
      .out(par_done_reg1502_out),
      .done(par_done_reg1502_done)
  );
  
  std_reg #(1) par_done_reg1503 (
      .in(par_done_reg1503_in),
      .write_en(par_done_reg1503_write_en),
      .clk(clk),
      .out(par_done_reg1503_out),
      .done(par_done_reg1503_done)
  );
  
  std_reg #(1) par_done_reg1504 (
      .in(par_done_reg1504_in),
      .write_en(par_done_reg1504_write_en),
      .clk(clk),
      .out(par_done_reg1504_out),
      .done(par_done_reg1504_done)
  );
  
  std_reg #(1) par_done_reg1505 (
      .in(par_done_reg1505_in),
      .write_en(par_done_reg1505_write_en),
      .clk(clk),
      .out(par_done_reg1505_out),
      .done(par_done_reg1505_done)
  );
  
  std_reg #(1) par_done_reg1506 (
      .in(par_done_reg1506_in),
      .write_en(par_done_reg1506_write_en),
      .clk(clk),
      .out(par_done_reg1506_out),
      .done(par_done_reg1506_done)
  );
  
  std_reg #(1) par_done_reg1507 (
      .in(par_done_reg1507_in),
      .write_en(par_done_reg1507_write_en),
      .clk(clk),
      .out(par_done_reg1507_out),
      .done(par_done_reg1507_done)
  );
  
  std_reg #(1) par_done_reg1508 (
      .in(par_done_reg1508_in),
      .write_en(par_done_reg1508_write_en),
      .clk(clk),
      .out(par_done_reg1508_out),
      .done(par_done_reg1508_done)
  );
  
  std_reg #(1) par_done_reg1509 (
      .in(par_done_reg1509_in),
      .write_en(par_done_reg1509_write_en),
      .clk(clk),
      .out(par_done_reg1509_out),
      .done(par_done_reg1509_done)
  );
  
  std_reg #(1) par_done_reg1510 (
      .in(par_done_reg1510_in),
      .write_en(par_done_reg1510_write_en),
      .clk(clk),
      .out(par_done_reg1510_out),
      .done(par_done_reg1510_done)
  );
  
  std_reg #(1) par_done_reg1511 (
      .in(par_done_reg1511_in),
      .write_en(par_done_reg1511_write_en),
      .clk(clk),
      .out(par_done_reg1511_out),
      .done(par_done_reg1511_done)
  );
  
  std_reg #(1) par_reset34 (
      .in(par_reset34_in),
      .write_en(par_reset34_write_en),
      .clk(clk),
      .out(par_reset34_out),
      .done(par_reset34_done)
  );
  
  std_reg #(1) par_done_reg1512 (
      .in(par_done_reg1512_in),
      .write_en(par_done_reg1512_write_en),
      .clk(clk),
      .out(par_done_reg1512_out),
      .done(par_done_reg1512_done)
  );
  
  std_reg #(1) par_done_reg1513 (
      .in(par_done_reg1513_in),
      .write_en(par_done_reg1513_write_en),
      .clk(clk),
      .out(par_done_reg1513_out),
      .done(par_done_reg1513_done)
  );
  
  std_reg #(1) par_done_reg1514 (
      .in(par_done_reg1514_in),
      .write_en(par_done_reg1514_write_en),
      .clk(clk),
      .out(par_done_reg1514_out),
      .done(par_done_reg1514_done)
  );
  
  std_reg #(1) par_done_reg1515 (
      .in(par_done_reg1515_in),
      .write_en(par_done_reg1515_write_en),
      .clk(clk),
      .out(par_done_reg1515_out),
      .done(par_done_reg1515_done)
  );
  
  std_reg #(1) par_done_reg1516 (
      .in(par_done_reg1516_in),
      .write_en(par_done_reg1516_write_en),
      .clk(clk),
      .out(par_done_reg1516_out),
      .done(par_done_reg1516_done)
  );
  
  std_reg #(1) par_done_reg1517 (
      .in(par_done_reg1517_in),
      .write_en(par_done_reg1517_write_en),
      .clk(clk),
      .out(par_done_reg1517_out),
      .done(par_done_reg1517_done)
  );
  
  std_reg #(1) par_done_reg1518 (
      .in(par_done_reg1518_in),
      .write_en(par_done_reg1518_write_en),
      .clk(clk),
      .out(par_done_reg1518_out),
      .done(par_done_reg1518_done)
  );
  
  std_reg #(1) par_done_reg1519 (
      .in(par_done_reg1519_in),
      .write_en(par_done_reg1519_write_en),
      .clk(clk),
      .out(par_done_reg1519_out),
      .done(par_done_reg1519_done)
  );
  
  std_reg #(1) par_done_reg1520 (
      .in(par_done_reg1520_in),
      .write_en(par_done_reg1520_write_en),
      .clk(clk),
      .out(par_done_reg1520_out),
      .done(par_done_reg1520_done)
  );
  
  std_reg #(1) par_done_reg1521 (
      .in(par_done_reg1521_in),
      .write_en(par_done_reg1521_write_en),
      .clk(clk),
      .out(par_done_reg1521_out),
      .done(par_done_reg1521_done)
  );
  
  std_reg #(1) par_done_reg1522 (
      .in(par_done_reg1522_in),
      .write_en(par_done_reg1522_write_en),
      .clk(clk),
      .out(par_done_reg1522_out),
      .done(par_done_reg1522_done)
  );
  
  std_reg #(1) par_done_reg1523 (
      .in(par_done_reg1523_in),
      .write_en(par_done_reg1523_write_en),
      .clk(clk),
      .out(par_done_reg1523_out),
      .done(par_done_reg1523_done)
  );
  
  std_reg #(1) par_done_reg1524 (
      .in(par_done_reg1524_in),
      .write_en(par_done_reg1524_write_en),
      .clk(clk),
      .out(par_done_reg1524_out),
      .done(par_done_reg1524_done)
  );
  
  std_reg #(1) par_done_reg1525 (
      .in(par_done_reg1525_in),
      .write_en(par_done_reg1525_write_en),
      .clk(clk),
      .out(par_done_reg1525_out),
      .done(par_done_reg1525_done)
  );
  
  std_reg #(1) par_done_reg1526 (
      .in(par_done_reg1526_in),
      .write_en(par_done_reg1526_write_en),
      .clk(clk),
      .out(par_done_reg1526_out),
      .done(par_done_reg1526_done)
  );
  
  std_reg #(1) par_done_reg1527 (
      .in(par_done_reg1527_in),
      .write_en(par_done_reg1527_write_en),
      .clk(clk),
      .out(par_done_reg1527_out),
      .done(par_done_reg1527_done)
  );
  
  std_reg #(1) par_done_reg1528 (
      .in(par_done_reg1528_in),
      .write_en(par_done_reg1528_write_en),
      .clk(clk),
      .out(par_done_reg1528_out),
      .done(par_done_reg1528_done)
  );
  
  std_reg #(1) par_done_reg1529 (
      .in(par_done_reg1529_in),
      .write_en(par_done_reg1529_write_en),
      .clk(clk),
      .out(par_done_reg1529_out),
      .done(par_done_reg1529_done)
  );
  
  std_reg #(1) par_done_reg1530 (
      .in(par_done_reg1530_in),
      .write_en(par_done_reg1530_write_en),
      .clk(clk),
      .out(par_done_reg1530_out),
      .done(par_done_reg1530_done)
  );
  
  std_reg #(1) par_done_reg1531 (
      .in(par_done_reg1531_in),
      .write_en(par_done_reg1531_write_en),
      .clk(clk),
      .out(par_done_reg1531_out),
      .done(par_done_reg1531_done)
  );
  
  std_reg #(1) par_done_reg1532 (
      .in(par_done_reg1532_in),
      .write_en(par_done_reg1532_write_en),
      .clk(clk),
      .out(par_done_reg1532_out),
      .done(par_done_reg1532_done)
  );
  
  std_reg #(1) par_done_reg1533 (
      .in(par_done_reg1533_in),
      .write_en(par_done_reg1533_write_en),
      .clk(clk),
      .out(par_done_reg1533_out),
      .done(par_done_reg1533_done)
  );
  
  std_reg #(1) par_done_reg1534 (
      .in(par_done_reg1534_in),
      .write_en(par_done_reg1534_write_en),
      .clk(clk),
      .out(par_done_reg1534_out),
      .done(par_done_reg1534_done)
  );
  
  std_reg #(1) par_done_reg1535 (
      .in(par_done_reg1535_in),
      .write_en(par_done_reg1535_write_en),
      .clk(clk),
      .out(par_done_reg1535_out),
      .done(par_done_reg1535_done)
  );
  
  std_reg #(1) par_done_reg1536 (
      .in(par_done_reg1536_in),
      .write_en(par_done_reg1536_write_en),
      .clk(clk),
      .out(par_done_reg1536_out),
      .done(par_done_reg1536_done)
  );
  
  std_reg #(1) par_done_reg1537 (
      .in(par_done_reg1537_in),
      .write_en(par_done_reg1537_write_en),
      .clk(clk),
      .out(par_done_reg1537_out),
      .done(par_done_reg1537_done)
  );
  
  std_reg #(1) par_done_reg1538 (
      .in(par_done_reg1538_in),
      .write_en(par_done_reg1538_write_en),
      .clk(clk),
      .out(par_done_reg1538_out),
      .done(par_done_reg1538_done)
  );
  
  std_reg #(1) par_done_reg1539 (
      .in(par_done_reg1539_in),
      .write_en(par_done_reg1539_write_en),
      .clk(clk),
      .out(par_done_reg1539_out),
      .done(par_done_reg1539_done)
  );
  
  std_reg #(1) par_done_reg1540 (
      .in(par_done_reg1540_in),
      .write_en(par_done_reg1540_write_en),
      .clk(clk),
      .out(par_done_reg1540_out),
      .done(par_done_reg1540_done)
  );
  
  std_reg #(1) par_done_reg1541 (
      .in(par_done_reg1541_in),
      .write_en(par_done_reg1541_write_en),
      .clk(clk),
      .out(par_done_reg1541_out),
      .done(par_done_reg1541_done)
  );
  
  std_reg #(1) par_done_reg1542 (
      .in(par_done_reg1542_in),
      .write_en(par_done_reg1542_write_en),
      .clk(clk),
      .out(par_done_reg1542_out),
      .done(par_done_reg1542_done)
  );
  
  std_reg #(1) par_done_reg1543 (
      .in(par_done_reg1543_in),
      .write_en(par_done_reg1543_write_en),
      .clk(clk),
      .out(par_done_reg1543_out),
      .done(par_done_reg1543_done)
  );
  
  std_reg #(1) par_done_reg1544 (
      .in(par_done_reg1544_in),
      .write_en(par_done_reg1544_write_en),
      .clk(clk),
      .out(par_done_reg1544_out),
      .done(par_done_reg1544_done)
  );
  
  std_reg #(1) par_done_reg1545 (
      .in(par_done_reg1545_in),
      .write_en(par_done_reg1545_write_en),
      .clk(clk),
      .out(par_done_reg1545_out),
      .done(par_done_reg1545_done)
  );
  
  std_reg #(1) par_done_reg1546 (
      .in(par_done_reg1546_in),
      .write_en(par_done_reg1546_write_en),
      .clk(clk),
      .out(par_done_reg1546_out),
      .done(par_done_reg1546_done)
  );
  
  std_reg #(1) par_done_reg1547 (
      .in(par_done_reg1547_in),
      .write_en(par_done_reg1547_write_en),
      .clk(clk),
      .out(par_done_reg1547_out),
      .done(par_done_reg1547_done)
  );
  
  std_reg #(1) par_done_reg1548 (
      .in(par_done_reg1548_in),
      .write_en(par_done_reg1548_write_en),
      .clk(clk),
      .out(par_done_reg1548_out),
      .done(par_done_reg1548_done)
  );
  
  std_reg #(1) par_done_reg1549 (
      .in(par_done_reg1549_in),
      .write_en(par_done_reg1549_write_en),
      .clk(clk),
      .out(par_done_reg1549_out),
      .done(par_done_reg1549_done)
  );
  
  std_reg #(1) par_done_reg1550 (
      .in(par_done_reg1550_in),
      .write_en(par_done_reg1550_write_en),
      .clk(clk),
      .out(par_done_reg1550_out),
      .done(par_done_reg1550_done)
  );
  
  std_reg #(1) par_done_reg1551 (
      .in(par_done_reg1551_in),
      .write_en(par_done_reg1551_write_en),
      .clk(clk),
      .out(par_done_reg1551_out),
      .done(par_done_reg1551_done)
  );
  
  std_reg #(1) par_done_reg1552 (
      .in(par_done_reg1552_in),
      .write_en(par_done_reg1552_write_en),
      .clk(clk),
      .out(par_done_reg1552_out),
      .done(par_done_reg1552_done)
  );
  
  std_reg #(1) par_done_reg1553 (
      .in(par_done_reg1553_in),
      .write_en(par_done_reg1553_write_en),
      .clk(clk),
      .out(par_done_reg1553_out),
      .done(par_done_reg1553_done)
  );
  
  std_reg #(1) par_reset35 (
      .in(par_reset35_in),
      .write_en(par_reset35_write_en),
      .clk(clk),
      .out(par_reset35_out),
      .done(par_reset35_done)
  );
  
  std_reg #(1) par_done_reg1554 (
      .in(par_done_reg1554_in),
      .write_en(par_done_reg1554_write_en),
      .clk(clk),
      .out(par_done_reg1554_out),
      .done(par_done_reg1554_done)
  );
  
  std_reg #(1) par_done_reg1555 (
      .in(par_done_reg1555_in),
      .write_en(par_done_reg1555_write_en),
      .clk(clk),
      .out(par_done_reg1555_out),
      .done(par_done_reg1555_done)
  );
  
  std_reg #(1) par_done_reg1556 (
      .in(par_done_reg1556_in),
      .write_en(par_done_reg1556_write_en),
      .clk(clk),
      .out(par_done_reg1556_out),
      .done(par_done_reg1556_done)
  );
  
  std_reg #(1) par_done_reg1557 (
      .in(par_done_reg1557_in),
      .write_en(par_done_reg1557_write_en),
      .clk(clk),
      .out(par_done_reg1557_out),
      .done(par_done_reg1557_done)
  );
  
  std_reg #(1) par_done_reg1558 (
      .in(par_done_reg1558_in),
      .write_en(par_done_reg1558_write_en),
      .clk(clk),
      .out(par_done_reg1558_out),
      .done(par_done_reg1558_done)
  );
  
  std_reg #(1) par_done_reg1559 (
      .in(par_done_reg1559_in),
      .write_en(par_done_reg1559_write_en),
      .clk(clk),
      .out(par_done_reg1559_out),
      .done(par_done_reg1559_done)
  );
  
  std_reg #(1) par_done_reg1560 (
      .in(par_done_reg1560_in),
      .write_en(par_done_reg1560_write_en),
      .clk(clk),
      .out(par_done_reg1560_out),
      .done(par_done_reg1560_done)
  );
  
  std_reg #(1) par_done_reg1561 (
      .in(par_done_reg1561_in),
      .write_en(par_done_reg1561_write_en),
      .clk(clk),
      .out(par_done_reg1561_out),
      .done(par_done_reg1561_done)
  );
  
  std_reg #(1) par_done_reg1562 (
      .in(par_done_reg1562_in),
      .write_en(par_done_reg1562_write_en),
      .clk(clk),
      .out(par_done_reg1562_out),
      .done(par_done_reg1562_done)
  );
  
  std_reg #(1) par_done_reg1563 (
      .in(par_done_reg1563_in),
      .write_en(par_done_reg1563_write_en),
      .clk(clk),
      .out(par_done_reg1563_out),
      .done(par_done_reg1563_done)
  );
  
  std_reg #(1) par_done_reg1564 (
      .in(par_done_reg1564_in),
      .write_en(par_done_reg1564_write_en),
      .clk(clk),
      .out(par_done_reg1564_out),
      .done(par_done_reg1564_done)
  );
  
  std_reg #(1) par_done_reg1565 (
      .in(par_done_reg1565_in),
      .write_en(par_done_reg1565_write_en),
      .clk(clk),
      .out(par_done_reg1565_out),
      .done(par_done_reg1565_done)
  );
  
  std_reg #(1) par_done_reg1566 (
      .in(par_done_reg1566_in),
      .write_en(par_done_reg1566_write_en),
      .clk(clk),
      .out(par_done_reg1566_out),
      .done(par_done_reg1566_done)
  );
  
  std_reg #(1) par_done_reg1567 (
      .in(par_done_reg1567_in),
      .write_en(par_done_reg1567_write_en),
      .clk(clk),
      .out(par_done_reg1567_out),
      .done(par_done_reg1567_done)
  );
  
  std_reg #(1) par_done_reg1568 (
      .in(par_done_reg1568_in),
      .write_en(par_done_reg1568_write_en),
      .clk(clk),
      .out(par_done_reg1568_out),
      .done(par_done_reg1568_done)
  );
  
  std_reg #(1) par_done_reg1569 (
      .in(par_done_reg1569_in),
      .write_en(par_done_reg1569_write_en),
      .clk(clk),
      .out(par_done_reg1569_out),
      .done(par_done_reg1569_done)
  );
  
  std_reg #(1) par_done_reg1570 (
      .in(par_done_reg1570_in),
      .write_en(par_done_reg1570_write_en),
      .clk(clk),
      .out(par_done_reg1570_out),
      .done(par_done_reg1570_done)
  );
  
  std_reg #(1) par_done_reg1571 (
      .in(par_done_reg1571_in),
      .write_en(par_done_reg1571_write_en),
      .clk(clk),
      .out(par_done_reg1571_out),
      .done(par_done_reg1571_done)
  );
  
  std_reg #(1) par_done_reg1572 (
      .in(par_done_reg1572_in),
      .write_en(par_done_reg1572_write_en),
      .clk(clk),
      .out(par_done_reg1572_out),
      .done(par_done_reg1572_done)
  );
  
  std_reg #(1) par_done_reg1573 (
      .in(par_done_reg1573_in),
      .write_en(par_done_reg1573_write_en),
      .clk(clk),
      .out(par_done_reg1573_out),
      .done(par_done_reg1573_done)
  );
  
  std_reg #(1) par_done_reg1574 (
      .in(par_done_reg1574_in),
      .write_en(par_done_reg1574_write_en),
      .clk(clk),
      .out(par_done_reg1574_out),
      .done(par_done_reg1574_done)
  );
  
  std_reg #(1) par_reset36 (
      .in(par_reset36_in),
      .write_en(par_reset36_write_en),
      .clk(clk),
      .out(par_reset36_out),
      .done(par_reset36_done)
  );
  
  std_reg #(1) par_done_reg1575 (
      .in(par_done_reg1575_in),
      .write_en(par_done_reg1575_write_en),
      .clk(clk),
      .out(par_done_reg1575_out),
      .done(par_done_reg1575_done)
  );
  
  std_reg #(1) par_done_reg1576 (
      .in(par_done_reg1576_in),
      .write_en(par_done_reg1576_write_en),
      .clk(clk),
      .out(par_done_reg1576_out),
      .done(par_done_reg1576_done)
  );
  
  std_reg #(1) par_done_reg1577 (
      .in(par_done_reg1577_in),
      .write_en(par_done_reg1577_write_en),
      .clk(clk),
      .out(par_done_reg1577_out),
      .done(par_done_reg1577_done)
  );
  
  std_reg #(1) par_done_reg1578 (
      .in(par_done_reg1578_in),
      .write_en(par_done_reg1578_write_en),
      .clk(clk),
      .out(par_done_reg1578_out),
      .done(par_done_reg1578_done)
  );
  
  std_reg #(1) par_done_reg1579 (
      .in(par_done_reg1579_in),
      .write_en(par_done_reg1579_write_en),
      .clk(clk),
      .out(par_done_reg1579_out),
      .done(par_done_reg1579_done)
  );
  
  std_reg #(1) par_done_reg1580 (
      .in(par_done_reg1580_in),
      .write_en(par_done_reg1580_write_en),
      .clk(clk),
      .out(par_done_reg1580_out),
      .done(par_done_reg1580_done)
  );
  
  std_reg #(1) par_done_reg1581 (
      .in(par_done_reg1581_in),
      .write_en(par_done_reg1581_write_en),
      .clk(clk),
      .out(par_done_reg1581_out),
      .done(par_done_reg1581_done)
  );
  
  std_reg #(1) par_done_reg1582 (
      .in(par_done_reg1582_in),
      .write_en(par_done_reg1582_write_en),
      .clk(clk),
      .out(par_done_reg1582_out),
      .done(par_done_reg1582_done)
  );
  
  std_reg #(1) par_done_reg1583 (
      .in(par_done_reg1583_in),
      .write_en(par_done_reg1583_write_en),
      .clk(clk),
      .out(par_done_reg1583_out),
      .done(par_done_reg1583_done)
  );
  
  std_reg #(1) par_done_reg1584 (
      .in(par_done_reg1584_in),
      .write_en(par_done_reg1584_write_en),
      .clk(clk),
      .out(par_done_reg1584_out),
      .done(par_done_reg1584_done)
  );
  
  std_reg #(1) par_done_reg1585 (
      .in(par_done_reg1585_in),
      .write_en(par_done_reg1585_write_en),
      .clk(clk),
      .out(par_done_reg1585_out),
      .done(par_done_reg1585_done)
  );
  
  std_reg #(1) par_done_reg1586 (
      .in(par_done_reg1586_in),
      .write_en(par_done_reg1586_write_en),
      .clk(clk),
      .out(par_done_reg1586_out),
      .done(par_done_reg1586_done)
  );
  
  std_reg #(1) par_done_reg1587 (
      .in(par_done_reg1587_in),
      .write_en(par_done_reg1587_write_en),
      .clk(clk),
      .out(par_done_reg1587_out),
      .done(par_done_reg1587_done)
  );
  
  std_reg #(1) par_done_reg1588 (
      .in(par_done_reg1588_in),
      .write_en(par_done_reg1588_write_en),
      .clk(clk),
      .out(par_done_reg1588_out),
      .done(par_done_reg1588_done)
  );
  
  std_reg #(1) par_done_reg1589 (
      .in(par_done_reg1589_in),
      .write_en(par_done_reg1589_write_en),
      .clk(clk),
      .out(par_done_reg1589_out),
      .done(par_done_reg1589_done)
  );
  
  std_reg #(1) par_done_reg1590 (
      .in(par_done_reg1590_in),
      .write_en(par_done_reg1590_write_en),
      .clk(clk),
      .out(par_done_reg1590_out),
      .done(par_done_reg1590_done)
  );
  
  std_reg #(1) par_done_reg1591 (
      .in(par_done_reg1591_in),
      .write_en(par_done_reg1591_write_en),
      .clk(clk),
      .out(par_done_reg1591_out),
      .done(par_done_reg1591_done)
  );
  
  std_reg #(1) par_done_reg1592 (
      .in(par_done_reg1592_in),
      .write_en(par_done_reg1592_write_en),
      .clk(clk),
      .out(par_done_reg1592_out),
      .done(par_done_reg1592_done)
  );
  
  std_reg #(1) par_done_reg1593 (
      .in(par_done_reg1593_in),
      .write_en(par_done_reg1593_write_en),
      .clk(clk),
      .out(par_done_reg1593_out),
      .done(par_done_reg1593_done)
  );
  
  std_reg #(1) par_done_reg1594 (
      .in(par_done_reg1594_in),
      .write_en(par_done_reg1594_write_en),
      .clk(clk),
      .out(par_done_reg1594_out),
      .done(par_done_reg1594_done)
  );
  
  std_reg #(1) par_done_reg1595 (
      .in(par_done_reg1595_in),
      .write_en(par_done_reg1595_write_en),
      .clk(clk),
      .out(par_done_reg1595_out),
      .done(par_done_reg1595_done)
  );
  
  std_reg #(1) par_done_reg1596 (
      .in(par_done_reg1596_in),
      .write_en(par_done_reg1596_write_en),
      .clk(clk),
      .out(par_done_reg1596_out),
      .done(par_done_reg1596_done)
  );
  
  std_reg #(1) par_done_reg1597 (
      .in(par_done_reg1597_in),
      .write_en(par_done_reg1597_write_en),
      .clk(clk),
      .out(par_done_reg1597_out),
      .done(par_done_reg1597_done)
  );
  
  std_reg #(1) par_done_reg1598 (
      .in(par_done_reg1598_in),
      .write_en(par_done_reg1598_write_en),
      .clk(clk),
      .out(par_done_reg1598_out),
      .done(par_done_reg1598_done)
  );
  
  std_reg #(1) par_done_reg1599 (
      .in(par_done_reg1599_in),
      .write_en(par_done_reg1599_write_en),
      .clk(clk),
      .out(par_done_reg1599_out),
      .done(par_done_reg1599_done)
  );
  
  std_reg #(1) par_done_reg1600 (
      .in(par_done_reg1600_in),
      .write_en(par_done_reg1600_write_en),
      .clk(clk),
      .out(par_done_reg1600_out),
      .done(par_done_reg1600_done)
  );
  
  std_reg #(1) par_done_reg1601 (
      .in(par_done_reg1601_in),
      .write_en(par_done_reg1601_write_en),
      .clk(clk),
      .out(par_done_reg1601_out),
      .done(par_done_reg1601_done)
  );
  
  std_reg #(1) par_done_reg1602 (
      .in(par_done_reg1602_in),
      .write_en(par_done_reg1602_write_en),
      .clk(clk),
      .out(par_done_reg1602_out),
      .done(par_done_reg1602_done)
  );
  
  std_reg #(1) par_done_reg1603 (
      .in(par_done_reg1603_in),
      .write_en(par_done_reg1603_write_en),
      .clk(clk),
      .out(par_done_reg1603_out),
      .done(par_done_reg1603_done)
  );
  
  std_reg #(1) par_done_reg1604 (
      .in(par_done_reg1604_in),
      .write_en(par_done_reg1604_write_en),
      .clk(clk),
      .out(par_done_reg1604_out),
      .done(par_done_reg1604_done)
  );
  
  std_reg #(1) par_reset37 (
      .in(par_reset37_in),
      .write_en(par_reset37_write_en),
      .clk(clk),
      .out(par_reset37_out),
      .done(par_reset37_done)
  );
  
  std_reg #(1) par_done_reg1605 (
      .in(par_done_reg1605_in),
      .write_en(par_done_reg1605_write_en),
      .clk(clk),
      .out(par_done_reg1605_out),
      .done(par_done_reg1605_done)
  );
  
  std_reg #(1) par_done_reg1606 (
      .in(par_done_reg1606_in),
      .write_en(par_done_reg1606_write_en),
      .clk(clk),
      .out(par_done_reg1606_out),
      .done(par_done_reg1606_done)
  );
  
  std_reg #(1) par_done_reg1607 (
      .in(par_done_reg1607_in),
      .write_en(par_done_reg1607_write_en),
      .clk(clk),
      .out(par_done_reg1607_out),
      .done(par_done_reg1607_done)
  );
  
  std_reg #(1) par_done_reg1608 (
      .in(par_done_reg1608_in),
      .write_en(par_done_reg1608_write_en),
      .clk(clk),
      .out(par_done_reg1608_out),
      .done(par_done_reg1608_done)
  );
  
  std_reg #(1) par_done_reg1609 (
      .in(par_done_reg1609_in),
      .write_en(par_done_reg1609_write_en),
      .clk(clk),
      .out(par_done_reg1609_out),
      .done(par_done_reg1609_done)
  );
  
  std_reg #(1) par_done_reg1610 (
      .in(par_done_reg1610_in),
      .write_en(par_done_reg1610_write_en),
      .clk(clk),
      .out(par_done_reg1610_out),
      .done(par_done_reg1610_done)
  );
  
  std_reg #(1) par_done_reg1611 (
      .in(par_done_reg1611_in),
      .write_en(par_done_reg1611_write_en),
      .clk(clk),
      .out(par_done_reg1611_out),
      .done(par_done_reg1611_done)
  );
  
  std_reg #(1) par_done_reg1612 (
      .in(par_done_reg1612_in),
      .write_en(par_done_reg1612_write_en),
      .clk(clk),
      .out(par_done_reg1612_out),
      .done(par_done_reg1612_done)
  );
  
  std_reg #(1) par_done_reg1613 (
      .in(par_done_reg1613_in),
      .write_en(par_done_reg1613_write_en),
      .clk(clk),
      .out(par_done_reg1613_out),
      .done(par_done_reg1613_done)
  );
  
  std_reg #(1) par_done_reg1614 (
      .in(par_done_reg1614_in),
      .write_en(par_done_reg1614_write_en),
      .clk(clk),
      .out(par_done_reg1614_out),
      .done(par_done_reg1614_done)
  );
  
  std_reg #(1) par_done_reg1615 (
      .in(par_done_reg1615_in),
      .write_en(par_done_reg1615_write_en),
      .clk(clk),
      .out(par_done_reg1615_out),
      .done(par_done_reg1615_done)
  );
  
  std_reg #(1) par_done_reg1616 (
      .in(par_done_reg1616_in),
      .write_en(par_done_reg1616_write_en),
      .clk(clk),
      .out(par_done_reg1616_out),
      .done(par_done_reg1616_done)
  );
  
  std_reg #(1) par_done_reg1617 (
      .in(par_done_reg1617_in),
      .write_en(par_done_reg1617_write_en),
      .clk(clk),
      .out(par_done_reg1617_out),
      .done(par_done_reg1617_done)
  );
  
  std_reg #(1) par_done_reg1618 (
      .in(par_done_reg1618_in),
      .write_en(par_done_reg1618_write_en),
      .clk(clk),
      .out(par_done_reg1618_out),
      .done(par_done_reg1618_done)
  );
  
  std_reg #(1) par_done_reg1619 (
      .in(par_done_reg1619_in),
      .write_en(par_done_reg1619_write_en),
      .clk(clk),
      .out(par_done_reg1619_out),
      .done(par_done_reg1619_done)
  );
  
  std_reg #(1) par_reset38 (
      .in(par_reset38_in),
      .write_en(par_reset38_write_en),
      .clk(clk),
      .out(par_reset38_out),
      .done(par_reset38_done)
  );
  
  std_reg #(1) par_done_reg1620 (
      .in(par_done_reg1620_in),
      .write_en(par_done_reg1620_write_en),
      .clk(clk),
      .out(par_done_reg1620_out),
      .done(par_done_reg1620_done)
  );
  
  std_reg #(1) par_done_reg1621 (
      .in(par_done_reg1621_in),
      .write_en(par_done_reg1621_write_en),
      .clk(clk),
      .out(par_done_reg1621_out),
      .done(par_done_reg1621_done)
  );
  
  std_reg #(1) par_done_reg1622 (
      .in(par_done_reg1622_in),
      .write_en(par_done_reg1622_write_en),
      .clk(clk),
      .out(par_done_reg1622_out),
      .done(par_done_reg1622_done)
  );
  
  std_reg #(1) par_done_reg1623 (
      .in(par_done_reg1623_in),
      .write_en(par_done_reg1623_write_en),
      .clk(clk),
      .out(par_done_reg1623_out),
      .done(par_done_reg1623_done)
  );
  
  std_reg #(1) par_done_reg1624 (
      .in(par_done_reg1624_in),
      .write_en(par_done_reg1624_write_en),
      .clk(clk),
      .out(par_done_reg1624_out),
      .done(par_done_reg1624_done)
  );
  
  std_reg #(1) par_done_reg1625 (
      .in(par_done_reg1625_in),
      .write_en(par_done_reg1625_write_en),
      .clk(clk),
      .out(par_done_reg1625_out),
      .done(par_done_reg1625_done)
  );
  
  std_reg #(1) par_done_reg1626 (
      .in(par_done_reg1626_in),
      .write_en(par_done_reg1626_write_en),
      .clk(clk),
      .out(par_done_reg1626_out),
      .done(par_done_reg1626_done)
  );
  
  std_reg #(1) par_done_reg1627 (
      .in(par_done_reg1627_in),
      .write_en(par_done_reg1627_write_en),
      .clk(clk),
      .out(par_done_reg1627_out),
      .done(par_done_reg1627_done)
  );
  
  std_reg #(1) par_done_reg1628 (
      .in(par_done_reg1628_in),
      .write_en(par_done_reg1628_write_en),
      .clk(clk),
      .out(par_done_reg1628_out),
      .done(par_done_reg1628_done)
  );
  
  std_reg #(1) par_done_reg1629 (
      .in(par_done_reg1629_in),
      .write_en(par_done_reg1629_write_en),
      .clk(clk),
      .out(par_done_reg1629_out),
      .done(par_done_reg1629_done)
  );
  
  std_reg #(1) par_done_reg1630 (
      .in(par_done_reg1630_in),
      .write_en(par_done_reg1630_write_en),
      .clk(clk),
      .out(par_done_reg1630_out),
      .done(par_done_reg1630_done)
  );
  
  std_reg #(1) par_done_reg1631 (
      .in(par_done_reg1631_in),
      .write_en(par_done_reg1631_write_en),
      .clk(clk),
      .out(par_done_reg1631_out),
      .done(par_done_reg1631_done)
  );
  
  std_reg #(1) par_done_reg1632 (
      .in(par_done_reg1632_in),
      .write_en(par_done_reg1632_write_en),
      .clk(clk),
      .out(par_done_reg1632_out),
      .done(par_done_reg1632_done)
  );
  
  std_reg #(1) par_done_reg1633 (
      .in(par_done_reg1633_in),
      .write_en(par_done_reg1633_write_en),
      .clk(clk),
      .out(par_done_reg1633_out),
      .done(par_done_reg1633_done)
  );
  
  std_reg #(1) par_done_reg1634 (
      .in(par_done_reg1634_in),
      .write_en(par_done_reg1634_write_en),
      .clk(clk),
      .out(par_done_reg1634_out),
      .done(par_done_reg1634_done)
  );
  
  std_reg #(1) par_done_reg1635 (
      .in(par_done_reg1635_in),
      .write_en(par_done_reg1635_write_en),
      .clk(clk),
      .out(par_done_reg1635_out),
      .done(par_done_reg1635_done)
  );
  
  std_reg #(1) par_done_reg1636 (
      .in(par_done_reg1636_in),
      .write_en(par_done_reg1636_write_en),
      .clk(clk),
      .out(par_done_reg1636_out),
      .done(par_done_reg1636_done)
  );
  
  std_reg #(1) par_done_reg1637 (
      .in(par_done_reg1637_in),
      .write_en(par_done_reg1637_write_en),
      .clk(clk),
      .out(par_done_reg1637_out),
      .done(par_done_reg1637_done)
  );
  
  std_reg #(1) par_done_reg1638 (
      .in(par_done_reg1638_in),
      .write_en(par_done_reg1638_write_en),
      .clk(clk),
      .out(par_done_reg1638_out),
      .done(par_done_reg1638_done)
  );
  
  std_reg #(1) par_done_reg1639 (
      .in(par_done_reg1639_in),
      .write_en(par_done_reg1639_write_en),
      .clk(clk),
      .out(par_done_reg1639_out),
      .done(par_done_reg1639_done)
  );
  
  std_reg #(1) par_reset39 (
      .in(par_reset39_in),
      .write_en(par_reset39_write_en),
      .clk(clk),
      .out(par_reset39_out),
      .done(par_reset39_done)
  );
  
  std_reg #(1) par_done_reg1640 (
      .in(par_done_reg1640_in),
      .write_en(par_done_reg1640_write_en),
      .clk(clk),
      .out(par_done_reg1640_out),
      .done(par_done_reg1640_done)
  );
  
  std_reg #(1) par_done_reg1641 (
      .in(par_done_reg1641_in),
      .write_en(par_done_reg1641_write_en),
      .clk(clk),
      .out(par_done_reg1641_out),
      .done(par_done_reg1641_done)
  );
  
  std_reg #(1) par_done_reg1642 (
      .in(par_done_reg1642_in),
      .write_en(par_done_reg1642_write_en),
      .clk(clk),
      .out(par_done_reg1642_out),
      .done(par_done_reg1642_done)
  );
  
  std_reg #(1) par_done_reg1643 (
      .in(par_done_reg1643_in),
      .write_en(par_done_reg1643_write_en),
      .clk(clk),
      .out(par_done_reg1643_out),
      .done(par_done_reg1643_done)
  );
  
  std_reg #(1) par_done_reg1644 (
      .in(par_done_reg1644_in),
      .write_en(par_done_reg1644_write_en),
      .clk(clk),
      .out(par_done_reg1644_out),
      .done(par_done_reg1644_done)
  );
  
  std_reg #(1) par_done_reg1645 (
      .in(par_done_reg1645_in),
      .write_en(par_done_reg1645_write_en),
      .clk(clk),
      .out(par_done_reg1645_out),
      .done(par_done_reg1645_done)
  );
  
  std_reg #(1) par_done_reg1646 (
      .in(par_done_reg1646_in),
      .write_en(par_done_reg1646_write_en),
      .clk(clk),
      .out(par_done_reg1646_out),
      .done(par_done_reg1646_done)
  );
  
  std_reg #(1) par_done_reg1647 (
      .in(par_done_reg1647_in),
      .write_en(par_done_reg1647_write_en),
      .clk(clk),
      .out(par_done_reg1647_out),
      .done(par_done_reg1647_done)
  );
  
  std_reg #(1) par_done_reg1648 (
      .in(par_done_reg1648_in),
      .write_en(par_done_reg1648_write_en),
      .clk(clk),
      .out(par_done_reg1648_out),
      .done(par_done_reg1648_done)
  );
  
  std_reg #(1) par_done_reg1649 (
      .in(par_done_reg1649_in),
      .write_en(par_done_reg1649_write_en),
      .clk(clk),
      .out(par_done_reg1649_out),
      .done(par_done_reg1649_done)
  );
  
  std_reg #(1) par_reset40 (
      .in(par_reset40_in),
      .write_en(par_reset40_write_en),
      .clk(clk),
      .out(par_reset40_out),
      .done(par_reset40_done)
  );
  
  std_reg #(1) par_done_reg1650 (
      .in(par_done_reg1650_in),
      .write_en(par_done_reg1650_write_en),
      .clk(clk),
      .out(par_done_reg1650_out),
      .done(par_done_reg1650_done)
  );
  
  std_reg #(1) par_done_reg1651 (
      .in(par_done_reg1651_in),
      .write_en(par_done_reg1651_write_en),
      .clk(clk),
      .out(par_done_reg1651_out),
      .done(par_done_reg1651_done)
  );
  
  std_reg #(1) par_done_reg1652 (
      .in(par_done_reg1652_in),
      .write_en(par_done_reg1652_write_en),
      .clk(clk),
      .out(par_done_reg1652_out),
      .done(par_done_reg1652_done)
  );
  
  std_reg #(1) par_done_reg1653 (
      .in(par_done_reg1653_in),
      .write_en(par_done_reg1653_write_en),
      .clk(clk),
      .out(par_done_reg1653_out),
      .done(par_done_reg1653_done)
  );
  
  std_reg #(1) par_done_reg1654 (
      .in(par_done_reg1654_in),
      .write_en(par_done_reg1654_write_en),
      .clk(clk),
      .out(par_done_reg1654_out),
      .done(par_done_reg1654_done)
  );
  
  std_reg #(1) par_done_reg1655 (
      .in(par_done_reg1655_in),
      .write_en(par_done_reg1655_write_en),
      .clk(clk),
      .out(par_done_reg1655_out),
      .done(par_done_reg1655_done)
  );
  
  std_reg #(1) par_done_reg1656 (
      .in(par_done_reg1656_in),
      .write_en(par_done_reg1656_write_en),
      .clk(clk),
      .out(par_done_reg1656_out),
      .done(par_done_reg1656_done)
  );
  
  std_reg #(1) par_done_reg1657 (
      .in(par_done_reg1657_in),
      .write_en(par_done_reg1657_write_en),
      .clk(clk),
      .out(par_done_reg1657_out),
      .done(par_done_reg1657_done)
  );
  
  std_reg #(1) par_done_reg1658 (
      .in(par_done_reg1658_in),
      .write_en(par_done_reg1658_write_en),
      .clk(clk),
      .out(par_done_reg1658_out),
      .done(par_done_reg1658_done)
  );
  
  std_reg #(1) par_done_reg1659 (
      .in(par_done_reg1659_in),
      .write_en(par_done_reg1659_write_en),
      .clk(clk),
      .out(par_done_reg1659_out),
      .done(par_done_reg1659_done)
  );
  
  std_reg #(1) par_done_reg1660 (
      .in(par_done_reg1660_in),
      .write_en(par_done_reg1660_write_en),
      .clk(clk),
      .out(par_done_reg1660_out),
      .done(par_done_reg1660_done)
  );
  
  std_reg #(1) par_done_reg1661 (
      .in(par_done_reg1661_in),
      .write_en(par_done_reg1661_write_en),
      .clk(clk),
      .out(par_done_reg1661_out),
      .done(par_done_reg1661_done)
  );
  
  std_reg #(1) par_reset41 (
      .in(par_reset41_in),
      .write_en(par_reset41_write_en),
      .clk(clk),
      .out(par_reset41_out),
      .done(par_reset41_done)
  );
  
  std_reg #(1) par_done_reg1662 (
      .in(par_done_reg1662_in),
      .write_en(par_done_reg1662_write_en),
      .clk(clk),
      .out(par_done_reg1662_out),
      .done(par_done_reg1662_done)
  );
  
  std_reg #(1) par_done_reg1663 (
      .in(par_done_reg1663_in),
      .write_en(par_done_reg1663_write_en),
      .clk(clk),
      .out(par_done_reg1663_out),
      .done(par_done_reg1663_done)
  );
  
  std_reg #(1) par_done_reg1664 (
      .in(par_done_reg1664_in),
      .write_en(par_done_reg1664_write_en),
      .clk(clk),
      .out(par_done_reg1664_out),
      .done(par_done_reg1664_done)
  );
  
  std_reg #(1) par_done_reg1665 (
      .in(par_done_reg1665_in),
      .write_en(par_done_reg1665_write_en),
      .clk(clk),
      .out(par_done_reg1665_out),
      .done(par_done_reg1665_done)
  );
  
  std_reg #(1) par_done_reg1666 (
      .in(par_done_reg1666_in),
      .write_en(par_done_reg1666_write_en),
      .clk(clk),
      .out(par_done_reg1666_out),
      .done(par_done_reg1666_done)
  );
  
  std_reg #(1) par_done_reg1667 (
      .in(par_done_reg1667_in),
      .write_en(par_done_reg1667_write_en),
      .clk(clk),
      .out(par_done_reg1667_out),
      .done(par_done_reg1667_done)
  );
  
  std_reg #(1) par_reset42 (
      .in(par_reset42_in),
      .write_en(par_reset42_write_en),
      .clk(clk),
      .out(par_reset42_out),
      .done(par_reset42_done)
  );
  
  std_reg #(1) par_done_reg1668 (
      .in(par_done_reg1668_in),
      .write_en(par_done_reg1668_write_en),
      .clk(clk),
      .out(par_done_reg1668_out),
      .done(par_done_reg1668_done)
  );
  
  std_reg #(1) par_done_reg1669 (
      .in(par_done_reg1669_in),
      .write_en(par_done_reg1669_write_en),
      .clk(clk),
      .out(par_done_reg1669_out),
      .done(par_done_reg1669_done)
  );
  
  std_reg #(1) par_done_reg1670 (
      .in(par_done_reg1670_in),
      .write_en(par_done_reg1670_write_en),
      .clk(clk),
      .out(par_done_reg1670_out),
      .done(par_done_reg1670_done)
  );
  
  std_reg #(1) par_done_reg1671 (
      .in(par_done_reg1671_in),
      .write_en(par_done_reg1671_write_en),
      .clk(clk),
      .out(par_done_reg1671_out),
      .done(par_done_reg1671_done)
  );
  
  std_reg #(1) par_done_reg1672 (
      .in(par_done_reg1672_in),
      .write_en(par_done_reg1672_write_en),
      .clk(clk),
      .out(par_done_reg1672_out),
      .done(par_done_reg1672_done)
  );
  
  std_reg #(1) par_done_reg1673 (
      .in(par_done_reg1673_in),
      .write_en(par_done_reg1673_write_en),
      .clk(clk),
      .out(par_done_reg1673_out),
      .done(par_done_reg1673_done)
  );
  
  std_reg #(1) par_reset43 (
      .in(par_reset43_in),
      .write_en(par_reset43_write_en),
      .clk(clk),
      .out(par_reset43_out),
      .done(par_reset43_done)
  );
  
  std_reg #(1) par_done_reg1674 (
      .in(par_done_reg1674_in),
      .write_en(par_done_reg1674_write_en),
      .clk(clk),
      .out(par_done_reg1674_out),
      .done(par_done_reg1674_done)
  );
  
  std_reg #(1) par_done_reg1675 (
      .in(par_done_reg1675_in),
      .write_en(par_done_reg1675_write_en),
      .clk(clk),
      .out(par_done_reg1675_out),
      .done(par_done_reg1675_done)
  );
  
  std_reg #(1) par_done_reg1676 (
      .in(par_done_reg1676_in),
      .write_en(par_done_reg1676_write_en),
      .clk(clk),
      .out(par_done_reg1676_out),
      .done(par_done_reg1676_done)
  );
  
  std_reg #(1) par_reset44 (
      .in(par_reset44_in),
      .write_en(par_reset44_write_en),
      .clk(clk),
      .out(par_reset44_out),
      .done(par_reset44_done)
  );
  
  std_reg #(1) par_done_reg1677 (
      .in(par_done_reg1677_in),
      .write_en(par_done_reg1677_write_en),
      .clk(clk),
      .out(par_done_reg1677_out),
      .done(par_done_reg1677_done)
  );
  
  std_reg #(1) par_done_reg1678 (
      .in(par_done_reg1678_in),
      .write_en(par_done_reg1678_write_en),
      .clk(clk),
      .out(par_done_reg1678_out),
      .done(par_done_reg1678_done)
  );
  
  std_reg #(1) par_reset45 (
      .in(par_reset45_in),
      .write_en(par_reset45_write_en),
      .clk(clk),
      .out(par_reset45_out),
      .done(par_reset45_done)
  );
  
  std_reg #(1) par_done_reg1679 (
      .in(par_done_reg1679_in),
      .write_en(par_done_reg1679_write_en),
      .clk(clk),
      .out(par_done_reg1679_out),
      .done(par_done_reg1679_done)
  );
  
  std_reg #(32) fsm0 (
      .in(fsm0_in),
      .write_en(fsm0_write_en),
      .clk(clk),
      .out(fsm0_out),
      .done(fsm0_done)
  );
  
  // Input / output connections
  assign done = (fsm0_out == 32'd110) ? 1'd1 : '0;
  assign out_mem_addr0 = (fsm0_out == 32'd102 & !out_mem_done & go | fsm0_out == 32'd103 & !out_mem_done & go | fsm0_out == 32'd104 & !out_mem_done & go | fsm0_out == 32'd105 & !out_mem_done & go | fsm0_out == 32'd106 & !out_mem_done & go | fsm0_out == 32'd107 & !out_mem_done & go | fsm0_out == 32'd108 & !out_mem_done & go | fsm0_out == 32'd109 & !out_mem_done & go) ? 4'd7 : (fsm0_out == 32'd94 & !out_mem_done & go | fsm0_out == 32'd95 & !out_mem_done & go | fsm0_out == 32'd96 & !out_mem_done & go | fsm0_out == 32'd97 & !out_mem_done & go | fsm0_out == 32'd98 & !out_mem_done & go | fsm0_out == 32'd99 & !out_mem_done & go | fsm0_out == 32'd100 & !out_mem_done & go | fsm0_out == 32'd101 & !out_mem_done & go) ? 4'd6 : (fsm0_out == 32'd86 & !out_mem_done & go | fsm0_out == 32'd87 & !out_mem_done & go | fsm0_out == 32'd88 & !out_mem_done & go | fsm0_out == 32'd89 & !out_mem_done & go | fsm0_out == 32'd90 & !out_mem_done & go | fsm0_out == 32'd91 & !out_mem_done & go | fsm0_out == 32'd92 & !out_mem_done & go | fsm0_out == 32'd93 & !out_mem_done & go) ? 4'd5 : (fsm0_out == 32'd78 & !out_mem_done & go | fsm0_out == 32'd79 & !out_mem_done & go | fsm0_out == 32'd80 & !out_mem_done & go | fsm0_out == 32'd81 & !out_mem_done & go | fsm0_out == 32'd82 & !out_mem_done & go | fsm0_out == 32'd83 & !out_mem_done & go | fsm0_out == 32'd84 & !out_mem_done & go | fsm0_out == 32'd85 & !out_mem_done & go) ? 4'd4 : (fsm0_out == 32'd70 & !out_mem_done & go | fsm0_out == 32'd71 & !out_mem_done & go | fsm0_out == 32'd72 & !out_mem_done & go | fsm0_out == 32'd73 & !out_mem_done & go | fsm0_out == 32'd74 & !out_mem_done & go | fsm0_out == 32'd75 & !out_mem_done & go | fsm0_out == 32'd76 & !out_mem_done & go | fsm0_out == 32'd77 & !out_mem_done & go) ? 4'd3 : (fsm0_out == 32'd62 & !out_mem_done & go | fsm0_out == 32'd63 & !out_mem_done & go | fsm0_out == 32'd64 & !out_mem_done & go | fsm0_out == 32'd65 & !out_mem_done & go | fsm0_out == 32'd66 & !out_mem_done & go | fsm0_out == 32'd67 & !out_mem_done & go | fsm0_out == 32'd68 & !out_mem_done & go | fsm0_out == 32'd69 & !out_mem_done & go) ? 4'd2 : (fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go | fsm0_out == 32'd53 & !out_mem_done & go) ? 4'd0 : (fsm0_out == 32'd54 & !out_mem_done & go | fsm0_out == 32'd55 & !out_mem_done & go | fsm0_out == 32'd56 & !out_mem_done & go | fsm0_out == 32'd57 & !out_mem_done & go | fsm0_out == 32'd58 & !out_mem_done & go | fsm0_out == 32'd59 & !out_mem_done & go | fsm0_out == 32'd60 & !out_mem_done & go | fsm0_out == 32'd61 & !out_mem_done & go) ? 4'd1 : '0;
  assign out_mem_addr1 = (fsm0_out == 32'd53 & !out_mem_done & go | fsm0_out == 32'd61 & !out_mem_done & go | fsm0_out == 32'd69 & !out_mem_done & go | fsm0_out == 32'd77 & !out_mem_done & go | fsm0_out == 32'd85 & !out_mem_done & go | fsm0_out == 32'd93 & !out_mem_done & go | fsm0_out == 32'd101 & !out_mem_done & go | fsm0_out == 32'd109 & !out_mem_done & go) ? 4'd7 : (fsm0_out == 32'd52 & !out_mem_done & go | fsm0_out == 32'd60 & !out_mem_done & go | fsm0_out == 32'd68 & !out_mem_done & go | fsm0_out == 32'd76 & !out_mem_done & go | fsm0_out == 32'd84 & !out_mem_done & go | fsm0_out == 32'd92 & !out_mem_done & go | fsm0_out == 32'd100 & !out_mem_done & go | fsm0_out == 32'd108 & !out_mem_done & go) ? 4'd6 : (fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd59 & !out_mem_done & go | fsm0_out == 32'd67 & !out_mem_done & go | fsm0_out == 32'd75 & !out_mem_done & go | fsm0_out == 32'd83 & !out_mem_done & go | fsm0_out == 32'd91 & !out_mem_done & go | fsm0_out == 32'd99 & !out_mem_done & go | fsm0_out == 32'd107 & !out_mem_done & go) ? 4'd5 : (fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd58 & !out_mem_done & go | fsm0_out == 32'd66 & !out_mem_done & go | fsm0_out == 32'd74 & !out_mem_done & go | fsm0_out == 32'd82 & !out_mem_done & go | fsm0_out == 32'd90 & !out_mem_done & go | fsm0_out == 32'd98 & !out_mem_done & go | fsm0_out == 32'd106 & !out_mem_done & go) ? 4'd4 : (fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd57 & !out_mem_done & go | fsm0_out == 32'd65 & !out_mem_done & go | fsm0_out == 32'd73 & !out_mem_done & go | fsm0_out == 32'd81 & !out_mem_done & go | fsm0_out == 32'd89 & !out_mem_done & go | fsm0_out == 32'd97 & !out_mem_done & go | fsm0_out == 32'd105 & !out_mem_done & go) ? 4'd3 : (fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd56 & !out_mem_done & go | fsm0_out == 32'd64 & !out_mem_done & go | fsm0_out == 32'd72 & !out_mem_done & go | fsm0_out == 32'd80 & !out_mem_done & go | fsm0_out == 32'd88 & !out_mem_done & go | fsm0_out == 32'd96 & !out_mem_done & go | fsm0_out == 32'd104 & !out_mem_done & go) ? 4'd2 : (fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd54 & !out_mem_done & go | fsm0_out == 32'd62 & !out_mem_done & go | fsm0_out == 32'd70 & !out_mem_done & go | fsm0_out == 32'd78 & !out_mem_done & go | fsm0_out == 32'd86 & !out_mem_done & go | fsm0_out == 32'd94 & !out_mem_done & go | fsm0_out == 32'd102 & !out_mem_done & go) ? 4'd0 : (fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd55 & !out_mem_done & go | fsm0_out == 32'd63 & !out_mem_done & go | fsm0_out == 32'd71 & !out_mem_done & go | fsm0_out == 32'd79 & !out_mem_done & go | fsm0_out == 32'd87 & !out_mem_done & go | fsm0_out == 32'd95 & !out_mem_done & go | fsm0_out == 32'd103 & !out_mem_done & go) ? 4'd1 : '0;
  assign out_mem_write_data = (fsm0_out == 32'd109 & !out_mem_done & go) ? pe_77_out : (fsm0_out == 32'd108 & !out_mem_done & go) ? pe_76_out : (fsm0_out == 32'd107 & !out_mem_done & go) ? pe_75_out : (fsm0_out == 32'd106 & !out_mem_done & go) ? pe_74_out : (fsm0_out == 32'd105 & !out_mem_done & go) ? pe_73_out : (fsm0_out == 32'd104 & !out_mem_done & go) ? pe_72_out : (fsm0_out == 32'd103 & !out_mem_done & go) ? pe_71_out : (fsm0_out == 32'd102 & !out_mem_done & go) ? pe_70_out : (fsm0_out == 32'd101 & !out_mem_done & go) ? pe_67_out : (fsm0_out == 32'd100 & !out_mem_done & go) ? pe_66_out : (fsm0_out == 32'd99 & !out_mem_done & go) ? pe_65_out : (fsm0_out == 32'd98 & !out_mem_done & go) ? pe_64_out : (fsm0_out == 32'd97 & !out_mem_done & go) ? pe_63_out : (fsm0_out == 32'd96 & !out_mem_done & go) ? pe_62_out : (fsm0_out == 32'd95 & !out_mem_done & go) ? pe_61_out : (fsm0_out == 32'd94 & !out_mem_done & go) ? pe_60_out : (fsm0_out == 32'd93 & !out_mem_done & go) ? pe_57_out : (fsm0_out == 32'd92 & !out_mem_done & go) ? pe_56_out : (fsm0_out == 32'd91 & !out_mem_done & go) ? pe_55_out : (fsm0_out == 32'd90 & !out_mem_done & go) ? pe_54_out : (fsm0_out == 32'd89 & !out_mem_done & go) ? pe_53_out : (fsm0_out == 32'd88 & !out_mem_done & go) ? pe_52_out : (fsm0_out == 32'd87 & !out_mem_done & go) ? pe_51_out : (fsm0_out == 32'd86 & !out_mem_done & go) ? pe_50_out : (fsm0_out == 32'd85 & !out_mem_done & go) ? pe_47_out : (fsm0_out == 32'd84 & !out_mem_done & go) ? pe_46_out : (fsm0_out == 32'd83 & !out_mem_done & go) ? pe_45_out : (fsm0_out == 32'd82 & !out_mem_done & go) ? pe_44_out : (fsm0_out == 32'd81 & !out_mem_done & go) ? pe_43_out : (fsm0_out == 32'd80 & !out_mem_done & go) ? pe_42_out : (fsm0_out == 32'd79 & !out_mem_done & go) ? pe_41_out : (fsm0_out == 32'd78 & !out_mem_done & go) ? pe_40_out : (fsm0_out == 32'd77 & !out_mem_done & go) ? pe_37_out : (fsm0_out == 32'd76 & !out_mem_done & go) ? pe_36_out : (fsm0_out == 32'd75 & !out_mem_done & go) ? pe_35_out : (fsm0_out == 32'd74 & !out_mem_done & go) ? pe_34_out : (fsm0_out == 32'd73 & !out_mem_done & go) ? pe_33_out : (fsm0_out == 32'd72 & !out_mem_done & go) ? pe_32_out : (fsm0_out == 32'd71 & !out_mem_done & go) ? pe_31_out : (fsm0_out == 32'd70 & !out_mem_done & go) ? pe_30_out : (fsm0_out == 32'd69 & !out_mem_done & go) ? pe_27_out : (fsm0_out == 32'd68 & !out_mem_done & go) ? pe_26_out : (fsm0_out == 32'd67 & !out_mem_done & go) ? pe_25_out : (fsm0_out == 32'd66 & !out_mem_done & go) ? pe_24_out : (fsm0_out == 32'd65 & !out_mem_done & go) ? pe_23_out : (fsm0_out == 32'd64 & !out_mem_done & go) ? pe_22_out : (fsm0_out == 32'd63 & !out_mem_done & go) ? pe_21_out : (fsm0_out == 32'd62 & !out_mem_done & go) ? pe_20_out : (fsm0_out == 32'd61 & !out_mem_done & go) ? pe_17_out : (fsm0_out == 32'd60 & !out_mem_done & go) ? pe_16_out : (fsm0_out == 32'd59 & !out_mem_done & go) ? pe_15_out : (fsm0_out == 32'd58 & !out_mem_done & go) ? pe_14_out : (fsm0_out == 32'd57 & !out_mem_done & go) ? pe_13_out : (fsm0_out == 32'd56 & !out_mem_done & go) ? pe_12_out : (fsm0_out == 32'd55 & !out_mem_done & go) ? pe_11_out : (fsm0_out == 32'd54 & !out_mem_done & go) ? pe_10_out : (fsm0_out == 32'd53 & !out_mem_done & go) ? pe_07_out : (fsm0_out == 32'd52 & !out_mem_done & go) ? pe_06_out : (fsm0_out == 32'd51 & !out_mem_done & go) ? pe_05_out : (fsm0_out == 32'd50 & !out_mem_done & go) ? pe_04_out : (fsm0_out == 32'd49 & !out_mem_done & go) ? pe_03_out : (fsm0_out == 32'd48 & !out_mem_done & go) ? pe_02_out : (fsm0_out == 32'd47 & !out_mem_done & go) ? pe_01_out : (fsm0_out == 32'd46 & !out_mem_done & go) ? pe_00_out : '0;
  assign out_mem_write_en = (fsm0_out == 32'd46 & !out_mem_done & go | fsm0_out == 32'd47 & !out_mem_done & go | fsm0_out == 32'd48 & !out_mem_done & go | fsm0_out == 32'd49 & !out_mem_done & go | fsm0_out == 32'd50 & !out_mem_done & go | fsm0_out == 32'd51 & !out_mem_done & go | fsm0_out == 32'd52 & !out_mem_done & go | fsm0_out == 32'd53 & !out_mem_done & go | fsm0_out == 32'd54 & !out_mem_done & go | fsm0_out == 32'd55 & !out_mem_done & go | fsm0_out == 32'd56 & !out_mem_done & go | fsm0_out == 32'd57 & !out_mem_done & go | fsm0_out == 32'd58 & !out_mem_done & go | fsm0_out == 32'd59 & !out_mem_done & go | fsm0_out == 32'd60 & !out_mem_done & go | fsm0_out == 32'd61 & !out_mem_done & go | fsm0_out == 32'd62 & !out_mem_done & go | fsm0_out == 32'd63 & !out_mem_done & go | fsm0_out == 32'd64 & !out_mem_done & go | fsm0_out == 32'd65 & !out_mem_done & go | fsm0_out == 32'd66 & !out_mem_done & go | fsm0_out == 32'd67 & !out_mem_done & go | fsm0_out == 32'd68 & !out_mem_done & go | fsm0_out == 32'd69 & !out_mem_done & go | fsm0_out == 32'd70 & !out_mem_done & go | fsm0_out == 32'd71 & !out_mem_done & go | fsm0_out == 32'd72 & !out_mem_done & go | fsm0_out == 32'd73 & !out_mem_done & go | fsm0_out == 32'd74 & !out_mem_done & go | fsm0_out == 32'd75 & !out_mem_done & go | fsm0_out == 32'd76 & !out_mem_done & go | fsm0_out == 32'd77 & !out_mem_done & go | fsm0_out == 32'd78 & !out_mem_done & go | fsm0_out == 32'd79 & !out_mem_done & go | fsm0_out == 32'd80 & !out_mem_done & go | fsm0_out == 32'd81 & !out_mem_done & go | fsm0_out == 32'd82 & !out_mem_done & go | fsm0_out == 32'd83 & !out_mem_done & go | fsm0_out == 32'd84 & !out_mem_done & go | fsm0_out == 32'd85 & !out_mem_done & go | fsm0_out == 32'd86 & !out_mem_done & go | fsm0_out == 32'd87 & !out_mem_done & go | fsm0_out == 32'd88 & !out_mem_done & go | fsm0_out == 32'd89 & !out_mem_done & go | fsm0_out == 32'd90 & !out_mem_done & go | fsm0_out == 32'd91 & !out_mem_done & go | fsm0_out == 32'd92 & !out_mem_done & go | fsm0_out == 32'd93 & !out_mem_done & go | fsm0_out == 32'd94 & !out_mem_done & go | fsm0_out == 32'd95 & !out_mem_done & go | fsm0_out == 32'd96 & !out_mem_done & go | fsm0_out == 32'd97 & !out_mem_done & go | fsm0_out == 32'd98 & !out_mem_done & go | fsm0_out == 32'd99 & !out_mem_done & go | fsm0_out == 32'd100 & !out_mem_done & go | fsm0_out == 32'd101 & !out_mem_done & go | fsm0_out == 32'd102 & !out_mem_done & go | fsm0_out == 32'd103 & !out_mem_done & go | fsm0_out == 32'd104 & !out_mem_done & go | fsm0_out == 32'd105 & !out_mem_done & go | fsm0_out == 32'd106 & !out_mem_done & go | fsm0_out == 32'd107 & !out_mem_done & go | fsm0_out == 32'd108 & !out_mem_done & go | fsm0_out == 32'd109 & !out_mem_done & go) ? 1'd1 : '0;
  assign left_77_read_in = (!(par_done_reg1391_out | left_77_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1483_out | left_77_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1553_out | left_77_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1604_out | left_77_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1639_out | left_77_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1661_out | left_77_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1673_out | left_77_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go | !(par_done_reg1678_out | left_77_read_done) & fsm0_out == 32'd44 & !par_reset44_out & go) ? right_76_write_out : '0;
  assign left_77_read_write_en = (!(par_done_reg1391_out | left_77_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1483_out | left_77_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1553_out | left_77_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1604_out | left_77_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1639_out | left_77_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1661_out | left_77_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1673_out | left_77_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go | !(par_done_reg1678_out | left_77_read_done) & fsm0_out == 32'd44 & !par_reset44_out & go) ? 1'd1 : '0;
  assign top_77_read_in = (!(par_done_reg1355_out | top_77_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1455_out | top_77_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1532_out | top_77_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1589_out | top_77_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1629_out | top_77_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1655_out | top_77_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1670_out | top_77_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go | !(par_done_reg1677_out | top_77_read_done) & fsm0_out == 32'd44 & !par_reset44_out & go) ? down_67_write_out : '0;
  assign top_77_read_write_en = (!(par_done_reg1355_out | top_77_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1455_out | top_77_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1532_out | top_77_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1589_out | top_77_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1629_out | top_77_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1655_out | top_77_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1670_out | top_77_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go | !(par_done_reg1677_out | top_77_read_done) & fsm0_out == 32'd44 & !par_reset44_out & go) ? 1'd1 : '0;
  assign pe_77_top = (!(par_done_reg1427_out | pe_77_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1511_out | pe_77_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1574_out | pe_77_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1619_out | pe_77_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1649_out | pe_77_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1667_out | pe_77_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1676_out | pe_77_done) & fsm0_out == 32'd43 & !par_reset43_out & go | !(par_done_reg1679_out | pe_77_done) & fsm0_out == 32'd45 & !par_reset45_out & go) ? top_77_read_out : '0;
  assign pe_77_left = (!(par_done_reg1427_out | pe_77_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1511_out | pe_77_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1574_out | pe_77_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1619_out | pe_77_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1649_out | pe_77_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1667_out | pe_77_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1676_out | pe_77_done) & fsm0_out == 32'd43 & !par_reset43_out & go | !(par_done_reg1679_out | pe_77_done) & fsm0_out == 32'd45 & !par_reset45_out & go) ? left_77_read_out : '0;
  assign pe_77_go = (!pe_77_done & (!(par_done_reg1427_out | pe_77_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1511_out | pe_77_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1574_out | pe_77_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1619_out | pe_77_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1649_out | pe_77_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1667_out | pe_77_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1676_out | pe_77_done) & fsm0_out == 32'd43 & !par_reset43_out & go | !(par_done_reg1679_out | pe_77_done) & fsm0_out == 32'd45 & !par_reset45_out & go)) ? 1'd1 : '0;
  assign right_76_write_in = (pe_76_done & (!(par_done_reg1319_out | right_76_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1426_out | right_76_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1510_out | right_76_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1573_out | right_76_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1618_out | right_76_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1648_out | right_76_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1666_out | right_76_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1675_out | right_76_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go)) ? pe_76_right : '0;
  assign right_76_write_write_en = (pe_76_done & (!(par_done_reg1319_out | right_76_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1426_out | right_76_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1510_out | right_76_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1573_out | right_76_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1618_out | right_76_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1648_out | right_76_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1666_out | right_76_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1675_out | right_76_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go)) ? 1'd1 : '0;
  assign left_76_read_in = (!(par_done_reg1275_out | left_76_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1390_out | left_76_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1482_out | left_76_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1552_out | left_76_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1603_out | left_76_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1638_out | left_76_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1660_out | left_76_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1672_out | left_76_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? right_75_write_out : '0;
  assign left_76_read_write_en = (!(par_done_reg1275_out | left_76_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1390_out | left_76_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1482_out | left_76_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1552_out | left_76_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1603_out | left_76_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1638_out | left_76_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1660_out | left_76_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1672_out | left_76_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign top_76_read_in = (!(par_done_reg1233_out | top_76_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1354_out | top_76_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1454_out | top_76_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1531_out | top_76_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1588_out | top_76_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1628_out | top_76_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1654_out | top_76_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1669_out | top_76_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? down_66_write_out : '0;
  assign top_76_read_write_en = (!(par_done_reg1233_out | top_76_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1354_out | top_76_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1454_out | top_76_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1531_out | top_76_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1588_out | top_76_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1628_out | top_76_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1654_out | top_76_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1669_out | top_76_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign pe_76_top = (!(par_done_reg1319_out | right_76_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1426_out | right_76_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1510_out | right_76_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1573_out | right_76_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1618_out | right_76_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1648_out | right_76_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1666_out | right_76_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1675_out | right_76_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go) ? top_76_read_out : '0;
  assign pe_76_left = (!(par_done_reg1319_out | right_76_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1426_out | right_76_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1510_out | right_76_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1573_out | right_76_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1618_out | right_76_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1648_out | right_76_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1666_out | right_76_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1675_out | right_76_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go) ? left_76_read_out : '0;
  assign pe_76_go = (!pe_76_done & (!(par_done_reg1319_out | right_76_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1426_out | right_76_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1510_out | right_76_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1573_out | right_76_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1618_out | right_76_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1648_out | right_76_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1666_out | right_76_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1675_out | right_76_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go)) ? 1'd1 : '0;
  assign right_75_write_in = (pe_75_done & (!(par_done_reg1191_out | right_75_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1318_out | right_75_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1425_out | right_75_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1509_out | right_75_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1572_out | right_75_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1617_out | right_75_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1647_out | right_75_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1665_out | right_75_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? pe_75_right : '0;
  assign right_75_write_write_en = (pe_75_done & (!(par_done_reg1191_out | right_75_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1318_out | right_75_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1425_out | right_75_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1509_out | right_75_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1572_out | right_75_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1617_out | right_75_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1647_out | right_75_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1665_out | right_75_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign left_75_read_in = (!(par_done_reg1141_out | left_75_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1274_out | left_75_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1389_out | left_75_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1481_out | left_75_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1551_out | left_75_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1602_out | left_75_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1637_out | left_75_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1659_out | left_75_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? right_74_write_out : '0;
  assign left_75_read_write_en = (!(par_done_reg1141_out | left_75_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1274_out | left_75_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1389_out | left_75_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1481_out | left_75_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1551_out | left_75_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1602_out | left_75_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1637_out | left_75_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1659_out | left_75_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign top_75_read_in = (!(par_done_reg1095_out | top_75_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1232_out | top_75_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1353_out | top_75_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1453_out | top_75_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1530_out | top_75_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1587_out | top_75_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1627_out | top_75_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1653_out | top_75_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? down_65_write_out : '0;
  assign top_75_read_write_en = (!(par_done_reg1095_out | top_75_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1232_out | top_75_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1353_out | top_75_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1453_out | top_75_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1530_out | top_75_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1587_out | top_75_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1627_out | top_75_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1653_out | top_75_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign pe_75_top = (!(par_done_reg1191_out | right_75_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1318_out | right_75_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1425_out | right_75_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1509_out | right_75_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1572_out | right_75_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1617_out | right_75_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1647_out | right_75_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1665_out | right_75_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go) ? top_75_read_out : '0;
  assign pe_75_left = (!(par_done_reg1191_out | right_75_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1318_out | right_75_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1425_out | right_75_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1509_out | right_75_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1572_out | right_75_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1617_out | right_75_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1647_out | right_75_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1665_out | right_75_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go) ? left_75_read_out : '0;
  assign pe_75_go = (!pe_75_done & (!(par_done_reg1191_out | right_75_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1318_out | right_75_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1425_out | right_75_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1509_out | right_75_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1572_out | right_75_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1617_out | right_75_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1647_out | right_75_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1665_out | right_75_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign right_74_write_in = (pe_74_done & (!(par_done_reg1049_out | right_74_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1190_out | right_74_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1317_out | right_74_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1424_out | right_74_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1508_out | right_74_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1571_out | right_74_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1616_out | right_74_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1646_out | right_74_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? pe_74_right : '0;
  assign right_74_write_write_en = (pe_74_done & (!(par_done_reg1049_out | right_74_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1190_out | right_74_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1317_out | right_74_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1424_out | right_74_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1508_out | right_74_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1571_out | right_74_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1616_out | right_74_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1646_out | right_74_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign left_74_read_in = (!(par_done_reg995_out | left_74_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1140_out | left_74_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1273_out | left_74_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1388_out | left_74_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1480_out | left_74_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1550_out | left_74_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1601_out | left_74_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1636_out | left_74_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? right_73_write_out : '0;
  assign left_74_read_write_en = (!(par_done_reg995_out | left_74_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1140_out | left_74_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1273_out | left_74_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1388_out | left_74_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1480_out | left_74_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1550_out | left_74_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1601_out | left_74_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1636_out | left_74_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign top_74_read_in = (!(par_done_reg947_out | top_74_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1094_out | top_74_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1231_out | top_74_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1352_out | top_74_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1452_out | top_74_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1529_out | top_74_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1586_out | top_74_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1626_out | top_74_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? down_64_write_out : '0;
  assign top_74_read_write_en = (!(par_done_reg947_out | top_74_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1094_out | top_74_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1231_out | top_74_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1352_out | top_74_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1452_out | top_74_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1529_out | top_74_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1586_out | top_74_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1626_out | top_74_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign pe_74_top = (!(par_done_reg1049_out | right_74_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1190_out | right_74_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1317_out | right_74_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1424_out | right_74_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1508_out | right_74_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1571_out | right_74_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1616_out | right_74_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1646_out | right_74_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? top_74_read_out : '0;
  assign pe_74_left = (!(par_done_reg1049_out | right_74_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1190_out | right_74_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1317_out | right_74_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1424_out | right_74_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1508_out | right_74_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1571_out | right_74_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1616_out | right_74_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1646_out | right_74_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? left_74_read_out : '0;
  assign pe_74_go = (!pe_74_done & (!(par_done_reg1049_out | right_74_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1190_out | right_74_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1317_out | right_74_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1424_out | right_74_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1508_out | right_74_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1571_out | right_74_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1616_out | right_74_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1646_out | right_74_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign right_73_write_in = (pe_73_done & (!(par_done_reg899_out | right_73_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1048_out | right_73_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1189_out | right_73_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1316_out | right_73_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1423_out | right_73_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1507_out | right_73_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1570_out | right_73_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1615_out | right_73_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_73_right : '0;
  assign right_73_write_write_en = (pe_73_done & (!(par_done_reg899_out | right_73_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1048_out | right_73_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1189_out | right_73_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1316_out | right_73_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1423_out | right_73_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1507_out | right_73_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1570_out | right_73_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1615_out | right_73_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign left_73_read_in = (!(par_done_reg843_out | left_73_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg994_out | left_73_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1139_out | left_73_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1272_out | left_73_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1387_out | left_73_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1479_out | left_73_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1549_out | left_73_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1600_out | left_73_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? right_72_write_out : '0;
  assign left_73_read_write_en = (!(par_done_reg843_out | left_73_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg994_out | left_73_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1139_out | left_73_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1272_out | left_73_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1387_out | left_73_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1479_out | left_73_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1549_out | left_73_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1600_out | left_73_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign top_73_read_in = (!(par_done_reg795_out | top_73_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg946_out | top_73_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1093_out | top_73_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1230_out | top_73_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1351_out | top_73_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1451_out | top_73_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1528_out | top_73_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1585_out | top_73_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? down_63_write_out : '0;
  assign top_73_read_write_en = (!(par_done_reg795_out | top_73_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg946_out | top_73_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1093_out | top_73_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1230_out | top_73_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1351_out | top_73_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1451_out | top_73_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1528_out | top_73_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1585_out | top_73_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign pe_73_top = (!(par_done_reg899_out | right_73_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1048_out | right_73_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1189_out | right_73_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1316_out | right_73_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1423_out | right_73_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1507_out | right_73_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1570_out | right_73_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1615_out | right_73_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? top_73_read_out : '0;
  assign pe_73_left = (!(par_done_reg899_out | right_73_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1048_out | right_73_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1189_out | right_73_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1316_out | right_73_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1423_out | right_73_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1507_out | right_73_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1570_out | right_73_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1615_out | right_73_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? left_73_read_out : '0;
  assign pe_73_go = (!pe_73_done & (!(par_done_reg899_out | right_73_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1048_out | right_73_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1189_out | right_73_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1316_out | right_73_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1423_out | right_73_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1507_out | right_73_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1570_out | right_73_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1615_out | right_73_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign right_72_write_in = (pe_72_done & (!(par_done_reg747_out | right_72_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg898_out | right_72_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1047_out | right_72_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1188_out | right_72_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1315_out | right_72_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1422_out | right_72_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1506_out | right_72_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1569_out | right_72_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_72_right : '0;
  assign right_72_write_write_en = (pe_72_done & (!(par_done_reg747_out | right_72_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg898_out | right_72_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1047_out | right_72_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1188_out | right_72_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1315_out | right_72_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1422_out | right_72_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1506_out | right_72_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1569_out | right_72_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign left_72_read_in = (!(par_done_reg691_out | left_72_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg842_out | left_72_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg993_out | left_72_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1138_out | left_72_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1271_out | left_72_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1386_out | left_72_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1478_out | left_72_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1548_out | left_72_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? right_71_write_out : '0;
  assign left_72_read_write_en = (!(par_done_reg691_out | left_72_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg842_out | left_72_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg993_out | left_72_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1138_out | left_72_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1271_out | left_72_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1386_out | left_72_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1478_out | left_72_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1548_out | left_72_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign top_72_read_in = (!(par_done_reg645_out | top_72_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg794_out | top_72_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg945_out | top_72_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1092_out | top_72_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1229_out | top_72_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1350_out | top_72_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1450_out | top_72_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1527_out | top_72_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? down_62_write_out : '0;
  assign top_72_read_write_en = (!(par_done_reg645_out | top_72_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg794_out | top_72_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg945_out | top_72_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1092_out | top_72_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1229_out | top_72_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1350_out | top_72_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1450_out | top_72_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1527_out | top_72_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign pe_72_top = (!(par_done_reg747_out | right_72_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg898_out | right_72_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1047_out | right_72_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1188_out | right_72_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1315_out | right_72_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1422_out | right_72_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1506_out | right_72_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1569_out | right_72_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? top_72_read_out : '0;
  assign pe_72_left = (!(par_done_reg747_out | right_72_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg898_out | right_72_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1047_out | right_72_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1188_out | right_72_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1315_out | right_72_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1422_out | right_72_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1506_out | right_72_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1569_out | right_72_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? left_72_read_out : '0;
  assign pe_72_go = (!pe_72_done & (!(par_done_reg747_out | right_72_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg898_out | right_72_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1047_out | right_72_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1188_out | right_72_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1315_out | right_72_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1422_out | right_72_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1506_out | right_72_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1569_out | right_72_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign right_71_write_in = (pe_71_done & (!(par_done_reg599_out | right_71_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg746_out | right_71_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg897_out | right_71_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1046_out | right_71_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1187_out | right_71_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1314_out | right_71_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1421_out | right_71_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1505_out | right_71_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_71_right : '0;
  assign right_71_write_write_en = (pe_71_done & (!(par_done_reg599_out | right_71_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg746_out | right_71_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg897_out | right_71_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1046_out | right_71_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1187_out | right_71_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1314_out | right_71_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1421_out | right_71_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1505_out | right_71_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_71_read_in = (!(par_done_reg545_out | left_71_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg690_out | left_71_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg841_out | left_71_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg992_out | left_71_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1137_out | left_71_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1270_out | left_71_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1385_out | left_71_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1477_out | left_71_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_70_write_out : '0;
  assign left_71_read_write_en = (!(par_done_reg545_out | left_71_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg690_out | left_71_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg841_out | left_71_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg992_out | left_71_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1137_out | left_71_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1270_out | left_71_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1385_out | left_71_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1477_out | left_71_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_71_read_in = (!(par_done_reg503_out | top_71_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg644_out | top_71_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg793_out | top_71_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg944_out | top_71_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1091_out | top_71_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1228_out | top_71_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1349_out | top_71_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1449_out | top_71_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_61_write_out : '0;
  assign top_71_read_write_en = (!(par_done_reg503_out | top_71_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg644_out | top_71_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg793_out | top_71_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg944_out | top_71_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1091_out | top_71_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1228_out | top_71_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1349_out | top_71_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1449_out | top_71_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_71_top = (!(par_done_reg599_out | right_71_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg746_out | right_71_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg897_out | right_71_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1046_out | right_71_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1187_out | right_71_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1314_out | right_71_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1421_out | right_71_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1505_out | right_71_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_71_read_out : '0;
  assign pe_71_left = (!(par_done_reg599_out | right_71_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg746_out | right_71_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg897_out | right_71_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1046_out | right_71_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1187_out | right_71_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1314_out | right_71_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1421_out | right_71_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1505_out | right_71_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_71_read_out : '0;
  assign pe_71_go = (!pe_71_done & (!(par_done_reg599_out | right_71_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg746_out | right_71_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg897_out | right_71_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1046_out | right_71_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1187_out | right_71_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1314_out | right_71_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1421_out | right_71_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1505_out | right_71_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_70_write_in = (pe_70_done & (!(par_done_reg461_out | right_70_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg598_out | right_70_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg745_out | right_70_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg896_out | right_70_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1045_out | right_70_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1186_out | right_70_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1313_out | right_70_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1420_out | right_70_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_70_right : '0;
  assign right_70_write_write_en = (pe_70_done & (!(par_done_reg461_out | right_70_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg598_out | right_70_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg745_out | right_70_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg896_out | right_70_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1045_out | right_70_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1186_out | right_70_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1313_out | right_70_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1420_out | right_70_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_70_read_in = (!(par_done_reg411_out | left_70_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg544_out | left_70_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg689_out | left_70_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg840_out | left_70_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg991_out | left_70_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1136_out | left_70_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1269_out | left_70_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1384_out | left_70_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? l7_read_data : '0;
  assign left_70_read_write_en = (!(par_done_reg411_out | left_70_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg544_out | left_70_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg689_out | left_70_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg840_out | left_70_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg991_out | left_70_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1136_out | left_70_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1269_out | left_70_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1384_out | left_70_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_70_read_in = (!(par_done_reg375_out | top_70_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg502_out | top_70_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg643_out | top_70_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg792_out | top_70_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg943_out | top_70_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1090_out | top_70_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1227_out | top_70_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1348_out | top_70_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_60_write_out : '0;
  assign top_70_read_write_en = (!(par_done_reg375_out | top_70_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg502_out | top_70_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg643_out | top_70_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg792_out | top_70_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg943_out | top_70_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1090_out | top_70_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1227_out | top_70_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1348_out | top_70_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_70_top = (!(par_done_reg461_out | right_70_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg598_out | right_70_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg745_out | right_70_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg896_out | right_70_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1045_out | right_70_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1186_out | right_70_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1313_out | right_70_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1420_out | right_70_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_70_read_out : '0;
  assign pe_70_left = (!(par_done_reg461_out | right_70_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg598_out | right_70_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg745_out | right_70_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg896_out | right_70_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1045_out | right_70_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1186_out | right_70_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1313_out | right_70_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1420_out | right_70_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_70_read_out : '0;
  assign pe_70_go = (!pe_70_done & (!(par_done_reg461_out | right_70_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg598_out | right_70_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg745_out | right_70_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg896_out | right_70_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1045_out | right_70_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1186_out | right_70_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1313_out | right_70_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1420_out | right_70_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_67_write_in = (pe_67_done & (!(par_done_reg1312_out | down_67_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1419_out | down_67_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1504_out | down_67_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1568_out | down_67_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1614_out | down_67_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1645_out | down_67_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1664_out | down_67_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1674_out | down_67_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go)) ? pe_67_down : '0;
  assign down_67_write_write_en = (pe_67_done & (!(par_done_reg1312_out | down_67_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1419_out | down_67_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1504_out | down_67_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1568_out | down_67_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1614_out | down_67_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1645_out | down_67_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1664_out | down_67_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1674_out | down_67_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go)) ? 1'd1 : '0;
  assign left_67_read_in = (!(par_done_reg1268_out | left_67_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1383_out | left_67_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1476_out | left_67_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1547_out | left_67_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1599_out | left_67_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1635_out | left_67_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1658_out | left_67_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1671_out | left_67_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? right_66_write_out : '0;
  assign left_67_read_write_en = (!(par_done_reg1268_out | left_67_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1383_out | left_67_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1476_out | left_67_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1547_out | left_67_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1599_out | left_67_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1635_out | left_67_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1658_out | left_67_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1671_out | left_67_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign top_67_read_in = (!(par_done_reg1226_out | top_67_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1347_out | top_67_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1448_out | top_67_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1526_out | top_67_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1584_out | top_67_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1625_out | top_67_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1652_out | top_67_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1668_out | top_67_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? down_57_write_out : '0;
  assign top_67_read_write_en = (!(par_done_reg1226_out | top_67_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1347_out | top_67_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1448_out | top_67_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1526_out | top_67_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1584_out | top_67_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1625_out | top_67_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1652_out | top_67_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go | !(par_done_reg1668_out | top_67_read_done) & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign pe_67_top = (!(par_done_reg1312_out | down_67_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1419_out | down_67_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1504_out | down_67_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1568_out | down_67_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1614_out | down_67_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1645_out | down_67_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1664_out | down_67_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1674_out | down_67_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go) ? top_67_read_out : '0;
  assign pe_67_left = (!(par_done_reg1312_out | down_67_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1419_out | down_67_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1504_out | down_67_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1568_out | down_67_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1614_out | down_67_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1645_out | down_67_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1664_out | down_67_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1674_out | down_67_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go) ? left_67_read_out : '0;
  assign pe_67_go = (!pe_67_done & (!(par_done_reg1312_out | down_67_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1419_out | down_67_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1504_out | down_67_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1568_out | down_67_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1614_out | down_67_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1645_out | down_67_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1664_out | down_67_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go | !(par_done_reg1674_out | down_67_write_done) & fsm0_out == 32'd43 & !par_reset43_out & go)) ? 1'd1 : '0;
  assign down_66_write_in = (pe_66_done & (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? pe_66_down : '0;
  assign down_66_write_write_en = (pe_66_done & (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign right_66_write_in = (pe_66_done & (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? pe_66_right : '0;
  assign right_66_write_write_en = (pe_66_done & (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign left_66_read_in = (!(par_done_reg1135_out | left_66_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1267_out | left_66_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1382_out | left_66_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1475_out | left_66_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1546_out | left_66_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1598_out | left_66_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1634_out | left_66_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1657_out | left_66_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? right_65_write_out : '0;
  assign left_66_read_write_en = (!(par_done_reg1135_out | left_66_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1267_out | left_66_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1382_out | left_66_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1475_out | left_66_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1546_out | left_66_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1598_out | left_66_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1634_out | left_66_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1657_out | left_66_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign top_66_read_in = (!(par_done_reg1089_out | top_66_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1225_out | top_66_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1346_out | top_66_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1447_out | top_66_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1525_out | top_66_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1583_out | top_66_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1624_out | top_66_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1651_out | top_66_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? down_56_write_out : '0;
  assign top_66_read_write_en = (!(par_done_reg1089_out | top_66_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1225_out | top_66_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1346_out | top_66_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1447_out | top_66_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1525_out | top_66_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1583_out | top_66_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1624_out | top_66_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1651_out | top_66_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign pe_66_top = (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go) ? top_66_read_out : '0;
  assign pe_66_left = (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go) ? left_66_read_out : '0;
  assign pe_66_go = (!pe_66_done & (!(par_done_reg1185_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1311_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1418_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1503_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1567_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1613_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1644_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1663_out | right_66_write_done & down_66_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign down_65_write_in = (pe_65_done & (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? pe_65_down : '0;
  assign down_65_write_write_en = (pe_65_done & (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign right_65_write_in = (pe_65_done & (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? pe_65_right : '0;
  assign right_65_write_write_en = (pe_65_done & (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign left_65_read_in = (!(par_done_reg990_out | left_65_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1134_out | left_65_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1266_out | left_65_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1381_out | left_65_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1474_out | left_65_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1545_out | left_65_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1597_out | left_65_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1633_out | left_65_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? right_64_write_out : '0;
  assign left_65_read_write_en = (!(par_done_reg990_out | left_65_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1134_out | left_65_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1266_out | left_65_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1381_out | left_65_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1474_out | left_65_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1545_out | left_65_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1597_out | left_65_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1633_out | left_65_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign top_65_read_in = (!(par_done_reg942_out | top_65_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1088_out | top_65_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1224_out | top_65_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1345_out | top_65_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1446_out | top_65_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1524_out | top_65_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1582_out | top_65_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1623_out | top_65_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? down_55_write_out : '0;
  assign top_65_read_write_en = (!(par_done_reg942_out | top_65_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1088_out | top_65_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1224_out | top_65_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1345_out | top_65_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1446_out | top_65_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1524_out | top_65_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1582_out | top_65_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1623_out | top_65_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign pe_65_top = (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? top_65_read_out : '0;
  assign pe_65_left = (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? left_65_read_out : '0;
  assign pe_65_go = (!pe_65_done & (!(par_done_reg1044_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1184_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1310_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1417_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1502_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1566_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1612_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1643_out | right_65_write_done & down_65_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign down_64_write_in = (pe_64_done & (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_64_down : '0;
  assign down_64_write_write_en = (pe_64_done & (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign right_64_write_in = (pe_64_done & (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_64_right : '0;
  assign right_64_write_write_en = (pe_64_done & (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign left_64_read_in = (!(par_done_reg839_out | left_64_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg989_out | left_64_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1133_out | left_64_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1265_out | left_64_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1380_out | left_64_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1473_out | left_64_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1544_out | left_64_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1596_out | left_64_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? right_63_write_out : '0;
  assign left_64_read_write_en = (!(par_done_reg839_out | left_64_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg989_out | left_64_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1133_out | left_64_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1265_out | left_64_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1380_out | left_64_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1473_out | left_64_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1544_out | left_64_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1596_out | left_64_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign top_64_read_in = (!(par_done_reg791_out | top_64_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg941_out | top_64_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1087_out | top_64_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1223_out | top_64_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1344_out | top_64_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1445_out | top_64_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1523_out | top_64_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1581_out | top_64_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? down_54_write_out : '0;
  assign top_64_read_write_en = (!(par_done_reg791_out | top_64_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg941_out | top_64_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1087_out | top_64_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1223_out | top_64_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1344_out | top_64_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1445_out | top_64_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1523_out | top_64_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1581_out | top_64_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign pe_64_top = (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? top_64_read_out : '0;
  assign pe_64_left = (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? left_64_read_out : '0;
  assign pe_64_go = (!pe_64_done & (!(par_done_reg895_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1043_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1183_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1309_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1416_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1501_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1565_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1611_out | right_64_write_done & down_64_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign down_63_write_in = (pe_63_done & (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_63_down : '0;
  assign down_63_write_write_en = (pe_63_done & (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign right_63_write_in = (pe_63_done & (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_63_right : '0;
  assign right_63_write_write_en = (pe_63_done & (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign left_63_read_in = (!(par_done_reg688_out | left_63_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg838_out | left_63_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg988_out | left_63_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1132_out | left_63_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1264_out | left_63_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1379_out | left_63_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1472_out | left_63_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1543_out | left_63_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? right_62_write_out : '0;
  assign left_63_read_write_en = (!(par_done_reg688_out | left_63_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg838_out | left_63_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg988_out | left_63_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1132_out | left_63_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1264_out | left_63_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1379_out | left_63_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1472_out | left_63_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1543_out | left_63_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign top_63_read_in = (!(par_done_reg642_out | top_63_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg790_out | top_63_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg940_out | top_63_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1086_out | top_63_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1222_out | top_63_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1343_out | top_63_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1444_out | top_63_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1522_out | top_63_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? down_53_write_out : '0;
  assign top_63_read_write_en = (!(par_done_reg642_out | top_63_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg790_out | top_63_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg940_out | top_63_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1086_out | top_63_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1222_out | top_63_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1343_out | top_63_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1444_out | top_63_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1522_out | top_63_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign pe_63_top = (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? top_63_read_out : '0;
  assign pe_63_left = (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? left_63_read_out : '0;
  assign pe_63_go = (!pe_63_done & (!(par_done_reg744_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg894_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1042_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1182_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1308_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1415_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1500_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1564_out | right_63_write_done & down_63_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign down_62_write_in = (pe_62_done & (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_62_down : '0;
  assign down_62_write_write_en = (pe_62_done & (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_62_write_in = (pe_62_done & (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_62_right : '0;
  assign right_62_write_write_en = (pe_62_done & (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_62_read_in = (!(par_done_reg543_out | left_62_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg687_out | left_62_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg837_out | left_62_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg987_out | left_62_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1131_out | left_62_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1263_out | left_62_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1378_out | left_62_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1471_out | left_62_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_61_write_out : '0;
  assign left_62_read_write_en = (!(par_done_reg543_out | left_62_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg687_out | left_62_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg837_out | left_62_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg987_out | left_62_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1131_out | left_62_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1263_out | left_62_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1378_out | left_62_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1471_out | left_62_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_62_read_in = (!(par_done_reg501_out | top_62_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg641_out | top_62_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg789_out | top_62_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg939_out | top_62_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1085_out | top_62_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1221_out | top_62_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1342_out | top_62_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1443_out | top_62_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_52_write_out : '0;
  assign top_62_read_write_en = (!(par_done_reg501_out | top_62_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg641_out | top_62_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg789_out | top_62_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg939_out | top_62_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1085_out | top_62_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1221_out | top_62_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1342_out | top_62_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1443_out | top_62_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_62_top = (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_62_read_out : '0;
  assign pe_62_left = (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_62_read_out : '0;
  assign pe_62_go = (!pe_62_done & (!(par_done_reg597_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg743_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg893_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1041_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1181_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1307_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1414_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1499_out | right_62_write_done & down_62_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign down_61_write_in = (pe_61_done & (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_61_down : '0;
  assign down_61_write_write_en = (pe_61_done & (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_61_write_in = (pe_61_done & (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_61_right : '0;
  assign right_61_write_write_en = (pe_61_done & (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_61_read_in = (!(par_done_reg410_out | left_61_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg542_out | left_61_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg686_out | left_61_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg836_out | left_61_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg986_out | left_61_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1130_out | left_61_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1262_out | left_61_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1377_out | left_61_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_60_write_out : '0;
  assign left_61_read_write_en = (!(par_done_reg410_out | left_61_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg542_out | left_61_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg686_out | left_61_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg836_out | left_61_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg986_out | left_61_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1130_out | left_61_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1262_out | left_61_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1377_out | left_61_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_61_read_in = (!(par_done_reg374_out | top_61_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg500_out | top_61_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg640_out | top_61_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg788_out | top_61_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg938_out | top_61_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1084_out | top_61_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1220_out | top_61_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1341_out | top_61_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_51_write_out : '0;
  assign top_61_read_write_en = (!(par_done_reg374_out | top_61_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg500_out | top_61_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg640_out | top_61_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg788_out | top_61_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg938_out | top_61_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1084_out | top_61_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1220_out | top_61_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1341_out | top_61_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_61_top = (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_61_read_out : '0;
  assign pe_61_left = (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_61_read_out : '0;
  assign pe_61_go = (!pe_61_done & (!(par_done_reg460_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg596_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg742_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg892_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1040_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1180_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1306_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1413_out | right_61_write_done & down_61_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_60_write_in = (pe_60_done & (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_60_down : '0;
  assign down_60_write_write_en = (pe_60_done & (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_60_write_in = (pe_60_done & (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_60_right : '0;
  assign right_60_write_write_en = (pe_60_done & (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_60_read_in = (!(par_done_reg295_out | left_60_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg409_out | left_60_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg541_out | left_60_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg685_out | left_60_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg835_out | left_60_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg985_out | left_60_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1129_out | left_60_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1261_out | left_60_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? l6_read_data : '0;
  assign left_60_read_write_en = (!(par_done_reg295_out | left_60_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg409_out | left_60_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg541_out | left_60_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg685_out | left_60_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg835_out | left_60_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg985_out | left_60_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1129_out | left_60_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1261_out | left_60_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_60_read_in = (!(par_done_reg267_out | top_60_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg373_out | top_60_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg499_out | top_60_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg639_out | top_60_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg787_out | top_60_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg937_out | top_60_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1083_out | top_60_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1219_out | top_60_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_50_write_out : '0;
  assign top_60_read_write_en = (!(par_done_reg267_out | top_60_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg373_out | top_60_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg499_out | top_60_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg639_out | top_60_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg787_out | top_60_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg937_out | top_60_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1083_out | top_60_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1219_out | top_60_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_60_top = (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_60_read_out : '0;
  assign pe_60_left = (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_60_read_out : '0;
  assign pe_60_go = (!pe_60_done & (!(par_done_reg339_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg459_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg595_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg741_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg891_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1039_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1179_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1305_out | right_60_write_done & down_60_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_57_write_in = (pe_57_done & (!(par_done_reg1178_out | down_57_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1304_out | down_57_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1412_out | down_57_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1498_out | down_57_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1563_out | down_57_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1610_out | down_57_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1642_out | down_57_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1662_out | down_57_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? pe_57_down : '0;
  assign down_57_write_write_en = (pe_57_done & (!(par_done_reg1178_out | down_57_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1304_out | down_57_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1412_out | down_57_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1498_out | down_57_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1563_out | down_57_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1610_out | down_57_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1642_out | down_57_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1662_out | down_57_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign left_57_read_in = (!(par_done_reg1128_out | left_57_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1260_out | left_57_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1376_out | left_57_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1470_out | left_57_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1542_out | left_57_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1595_out | left_57_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1632_out | left_57_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1656_out | left_57_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? right_56_write_out : '0;
  assign left_57_read_write_en = (!(par_done_reg1128_out | left_57_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1260_out | left_57_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1376_out | left_57_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1470_out | left_57_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1542_out | left_57_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1595_out | left_57_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1632_out | left_57_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1656_out | left_57_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign top_57_read_in = (!(par_done_reg1082_out | top_57_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1218_out | top_57_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1340_out | top_57_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1442_out | top_57_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1521_out | top_57_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1580_out | top_57_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1622_out | top_57_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1650_out | top_57_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? down_47_write_out : '0;
  assign top_57_read_write_en = (!(par_done_reg1082_out | top_57_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1218_out | top_57_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1340_out | top_57_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1442_out | top_57_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1521_out | top_57_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1580_out | top_57_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1622_out | top_57_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go | !(par_done_reg1650_out | top_57_read_done) & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign pe_57_top = (!(par_done_reg1178_out | down_57_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1304_out | down_57_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1412_out | down_57_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1498_out | down_57_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1563_out | down_57_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1610_out | down_57_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1642_out | down_57_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1662_out | down_57_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go) ? top_57_read_out : '0;
  assign pe_57_left = (!(par_done_reg1178_out | down_57_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1304_out | down_57_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1412_out | down_57_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1498_out | down_57_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1563_out | down_57_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1610_out | down_57_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1642_out | down_57_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1662_out | down_57_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go) ? left_57_read_out : '0;
  assign pe_57_go = (!pe_57_done & (!(par_done_reg1178_out | down_57_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1304_out | down_57_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1412_out | down_57_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1498_out | down_57_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1563_out | down_57_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1610_out | down_57_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1642_out | down_57_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go | !(par_done_reg1662_out | down_57_write_done) & fsm0_out == 32'd41 & !par_reset41_out & go)) ? 1'd1 : '0;
  assign down_56_write_in = (pe_56_done & (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? pe_56_down : '0;
  assign down_56_write_write_en = (pe_56_done & (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign right_56_write_in = (pe_56_done & (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? pe_56_right : '0;
  assign right_56_write_write_en = (pe_56_done & (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign left_56_read_in = (!(par_done_reg984_out | left_56_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1127_out | left_56_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1259_out | left_56_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1375_out | left_56_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1469_out | left_56_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1541_out | left_56_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1594_out | left_56_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1631_out | left_56_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? right_55_write_out : '0;
  assign left_56_read_write_en = (!(par_done_reg984_out | left_56_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1127_out | left_56_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1259_out | left_56_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1375_out | left_56_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1469_out | left_56_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1541_out | left_56_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1594_out | left_56_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1631_out | left_56_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign top_56_read_in = (!(par_done_reg936_out | top_56_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1081_out | top_56_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1217_out | top_56_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1339_out | top_56_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1441_out | top_56_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1520_out | top_56_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1579_out | top_56_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1621_out | top_56_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? down_46_write_out : '0;
  assign top_56_read_write_en = (!(par_done_reg936_out | top_56_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1081_out | top_56_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1217_out | top_56_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1339_out | top_56_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1441_out | top_56_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1520_out | top_56_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1579_out | top_56_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1621_out | top_56_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign pe_56_top = (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? top_56_read_out : '0;
  assign pe_56_left = (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? left_56_read_out : '0;
  assign pe_56_go = (!pe_56_done & (!(par_done_reg1038_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1177_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1303_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1411_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1497_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1562_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1609_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1641_out | right_56_write_done & down_56_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign down_55_write_in = (pe_55_done & (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_55_down : '0;
  assign down_55_write_write_en = (pe_55_done & (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign right_55_write_in = (pe_55_done & (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_55_right : '0;
  assign right_55_write_write_en = (pe_55_done & (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign left_55_read_in = (!(par_done_reg834_out | left_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg983_out | left_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1126_out | left_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1258_out | left_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1374_out | left_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1468_out | left_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1540_out | left_55_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1593_out | left_55_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? right_54_write_out : '0;
  assign left_55_read_write_en = (!(par_done_reg834_out | left_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg983_out | left_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1126_out | left_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1258_out | left_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1374_out | left_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1468_out | left_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1540_out | left_55_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1593_out | left_55_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign top_55_read_in = (!(par_done_reg786_out | top_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg935_out | top_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1080_out | top_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1216_out | top_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1338_out | top_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1440_out | top_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1519_out | top_55_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1578_out | top_55_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? down_45_write_out : '0;
  assign top_55_read_write_en = (!(par_done_reg786_out | top_55_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg935_out | top_55_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1080_out | top_55_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1216_out | top_55_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1338_out | top_55_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1440_out | top_55_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1519_out | top_55_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1578_out | top_55_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign pe_55_top = (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? top_55_read_out : '0;
  assign pe_55_left = (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? left_55_read_out : '0;
  assign pe_55_go = (!pe_55_done & (!(par_done_reg890_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1037_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1176_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1302_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1410_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1496_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1561_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1608_out | right_55_write_done & down_55_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign down_54_write_in = (pe_54_done & (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_54_down : '0;
  assign down_54_write_write_en = (pe_54_done & (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign right_54_write_in = (pe_54_done & (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_54_right : '0;
  assign right_54_write_write_en = (pe_54_done & (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign left_54_read_in = (!(par_done_reg684_out | left_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg833_out | left_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg982_out | left_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1125_out | left_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1257_out | left_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1373_out | left_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1467_out | left_54_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1539_out | left_54_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? right_53_write_out : '0;
  assign left_54_read_write_en = (!(par_done_reg684_out | left_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg833_out | left_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg982_out | left_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1125_out | left_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1257_out | left_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1373_out | left_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1467_out | left_54_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1539_out | left_54_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign top_54_read_in = (!(par_done_reg638_out | top_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg785_out | top_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg934_out | top_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1079_out | top_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1215_out | top_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1337_out | top_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1439_out | top_54_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1518_out | top_54_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? down_44_write_out : '0;
  assign top_54_read_write_en = (!(par_done_reg638_out | top_54_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg785_out | top_54_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg934_out | top_54_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1079_out | top_54_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1215_out | top_54_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1337_out | top_54_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1439_out | top_54_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1518_out | top_54_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign pe_54_top = (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? top_54_read_out : '0;
  assign pe_54_left = (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? left_54_read_out : '0;
  assign pe_54_go = (!pe_54_done & (!(par_done_reg740_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg889_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1036_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1175_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1301_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1409_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1495_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1560_out | right_54_write_done & down_54_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign down_53_write_in = (pe_53_done & (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_53_down : '0;
  assign down_53_write_write_en = (pe_53_done & (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_53_write_in = (pe_53_done & (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_53_right : '0;
  assign right_53_write_write_en = (pe_53_done & (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_53_read_in = (!(par_done_reg540_out | left_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg683_out | left_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg832_out | left_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg981_out | left_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1124_out | left_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1256_out | left_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1372_out | left_53_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1466_out | left_53_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_52_write_out : '0;
  assign left_53_read_write_en = (!(par_done_reg540_out | left_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg683_out | left_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg832_out | left_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg981_out | left_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1124_out | left_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1256_out | left_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1372_out | left_53_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1466_out | left_53_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_53_read_in = (!(par_done_reg498_out | top_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg637_out | top_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg784_out | top_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg933_out | top_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1078_out | top_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1214_out | top_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1336_out | top_53_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1438_out | top_53_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_43_write_out : '0;
  assign top_53_read_write_en = (!(par_done_reg498_out | top_53_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg637_out | top_53_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg784_out | top_53_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg933_out | top_53_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1078_out | top_53_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1214_out | top_53_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1336_out | top_53_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1438_out | top_53_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_53_top = (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_53_read_out : '0;
  assign pe_53_left = (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_53_read_out : '0;
  assign pe_53_go = (!pe_53_done & (!(par_done_reg594_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg739_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg888_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1035_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1174_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1300_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1408_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1494_out | right_53_write_done & down_53_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign down_52_write_in = (pe_52_done & (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_52_down : '0;
  assign down_52_write_write_en = (pe_52_done & (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_52_write_in = (pe_52_done & (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_52_right : '0;
  assign right_52_write_write_en = (pe_52_done & (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_52_read_in = (!(par_done_reg408_out | left_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg539_out | left_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg682_out | left_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg831_out | left_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg980_out | left_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1123_out | left_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1255_out | left_52_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1371_out | left_52_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_51_write_out : '0;
  assign left_52_read_write_en = (!(par_done_reg408_out | left_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg539_out | left_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg682_out | left_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg831_out | left_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg980_out | left_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1123_out | left_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1255_out | left_52_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1371_out | left_52_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_52_read_in = (!(par_done_reg372_out | top_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg497_out | top_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg636_out | top_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg783_out | top_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg932_out | top_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1077_out | top_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1213_out | top_52_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1335_out | top_52_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_42_write_out : '0;
  assign top_52_read_write_en = (!(par_done_reg372_out | top_52_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg497_out | top_52_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg636_out | top_52_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg783_out | top_52_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg932_out | top_52_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1077_out | top_52_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1213_out | top_52_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1335_out | top_52_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_52_top = (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_52_read_out : '0;
  assign pe_52_left = (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_52_read_out : '0;
  assign pe_52_go = (!pe_52_done & (!(par_done_reg458_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg593_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg738_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg887_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1034_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1173_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1299_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1407_out | right_52_write_done & down_52_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_51_write_in = (pe_51_done & (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_51_down : '0;
  assign down_51_write_write_en = (pe_51_done & (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_51_write_in = (pe_51_done & (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_51_right : '0;
  assign right_51_write_write_en = (pe_51_done & (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_51_read_in = (!(par_done_reg294_out | left_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg407_out | left_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg538_out | left_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg681_out | left_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg830_out | left_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg979_out | left_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1122_out | left_51_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1254_out | left_51_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_50_write_out : '0;
  assign left_51_read_write_en = (!(par_done_reg294_out | left_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg407_out | left_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg538_out | left_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg681_out | left_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg830_out | left_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg979_out | left_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1122_out | left_51_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1254_out | left_51_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_51_read_in = (!(par_done_reg266_out | top_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg371_out | top_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg496_out | top_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg635_out | top_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg782_out | top_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg931_out | top_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1076_out | top_51_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1212_out | top_51_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_41_write_out : '0;
  assign top_51_read_write_en = (!(par_done_reg266_out | top_51_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg371_out | top_51_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg496_out | top_51_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg635_out | top_51_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg782_out | top_51_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg931_out | top_51_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1076_out | top_51_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1212_out | top_51_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_51_top = (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_51_read_out : '0;
  assign pe_51_left = (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_51_read_out : '0;
  assign pe_51_go = (!pe_51_done & (!(par_done_reg338_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg457_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg592_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg737_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg886_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1033_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1172_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1298_out | right_51_write_done & down_51_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_50_write_in = (pe_50_done & (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_50_down : '0;
  assign down_50_write_write_en = (pe_50_done & (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_50_write_in = (pe_50_done & (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_50_right : '0;
  assign right_50_write_write_en = (pe_50_done & (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_50_read_in = (!(par_done_reg204_out | left_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg293_out | left_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg406_out | left_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg537_out | left_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg680_out | left_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg829_out | left_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg978_out | left_50_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1121_out | left_50_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? l5_read_data : '0;
  assign left_50_read_write_en = (!(par_done_reg204_out | left_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg293_out | left_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg406_out | left_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg537_out | left_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg680_out | left_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg829_out | left_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg978_out | left_50_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1121_out | left_50_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_50_read_in = (!(par_done_reg183_out | top_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg265_out | top_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg370_out | top_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg495_out | top_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg634_out | top_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg781_out | top_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg930_out | top_50_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1075_out | top_50_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_40_write_out : '0;
  assign top_50_read_write_en = (!(par_done_reg183_out | top_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg265_out | top_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg370_out | top_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg495_out | top_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg634_out | top_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg781_out | top_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg930_out | top_50_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1075_out | top_50_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_50_top = (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_50_read_out : '0;
  assign pe_50_left = (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_50_read_out : '0;
  assign pe_50_go = (!pe_50_done & (!(par_done_reg239_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg337_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg456_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg591_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg736_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg885_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1032_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1171_out | right_50_write_done & down_50_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_47_write_in = (pe_47_done & (!(par_done_reg1031_out | down_47_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1170_out | down_47_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1297_out | down_47_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1406_out | down_47_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1493_out | down_47_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1559_out | down_47_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1607_out | down_47_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1640_out | down_47_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? pe_47_down : '0;
  assign down_47_write_write_en = (pe_47_done & (!(par_done_reg1031_out | down_47_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1170_out | down_47_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1297_out | down_47_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1406_out | down_47_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1493_out | down_47_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1559_out | down_47_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1607_out | down_47_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1640_out | down_47_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign left_47_read_in = (!(par_done_reg977_out | left_47_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1120_out | left_47_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1253_out | left_47_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1370_out | left_47_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1465_out | left_47_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1538_out | left_47_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1592_out | left_47_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1630_out | left_47_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? right_46_write_out : '0;
  assign left_47_read_write_en = (!(par_done_reg977_out | left_47_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1120_out | left_47_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1253_out | left_47_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1370_out | left_47_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1465_out | left_47_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1538_out | left_47_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1592_out | left_47_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1630_out | left_47_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign top_47_read_in = (!(par_done_reg929_out | top_47_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1074_out | top_47_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1211_out | top_47_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1334_out | top_47_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1437_out | top_47_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1517_out | top_47_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1577_out | top_47_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1620_out | top_47_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? down_37_write_out : '0;
  assign top_47_read_write_en = (!(par_done_reg929_out | top_47_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1074_out | top_47_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1211_out | top_47_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1334_out | top_47_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1437_out | top_47_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1517_out | top_47_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1577_out | top_47_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go | !(par_done_reg1620_out | top_47_read_done) & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign pe_47_top = (!(par_done_reg1031_out | down_47_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1170_out | down_47_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1297_out | down_47_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1406_out | down_47_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1493_out | down_47_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1559_out | down_47_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1607_out | down_47_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1640_out | down_47_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? top_47_read_out : '0;
  assign pe_47_left = (!(par_done_reg1031_out | down_47_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1170_out | down_47_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1297_out | down_47_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1406_out | down_47_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1493_out | down_47_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1559_out | down_47_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1607_out | down_47_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1640_out | down_47_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go) ? left_47_read_out : '0;
  assign pe_47_go = (!pe_47_done & (!(par_done_reg1031_out | down_47_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1170_out | down_47_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1297_out | down_47_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1406_out | down_47_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1493_out | down_47_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1559_out | down_47_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1607_out | down_47_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go | !(par_done_reg1640_out | down_47_write_done) & fsm0_out == 32'd39 & !par_reset39_out & go)) ? 1'd1 : '0;
  assign down_46_write_in = (pe_46_done & (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_46_down : '0;
  assign down_46_write_write_en = (pe_46_done & (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign right_46_write_in = (pe_46_done & (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_46_right : '0;
  assign right_46_write_write_en = (pe_46_done & (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign left_46_read_in = (!(par_done_reg828_out | left_46_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg976_out | left_46_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1119_out | left_46_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1252_out | left_46_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1369_out | left_46_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1464_out | left_46_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1537_out | left_46_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1591_out | left_46_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? right_45_write_out : '0;
  assign left_46_read_write_en = (!(par_done_reg828_out | left_46_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg976_out | left_46_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1119_out | left_46_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1252_out | left_46_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1369_out | left_46_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1464_out | left_46_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1537_out | left_46_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1591_out | left_46_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign top_46_read_in = (!(par_done_reg780_out | top_46_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg928_out | top_46_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1073_out | top_46_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1210_out | top_46_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1333_out | top_46_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1436_out | top_46_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1516_out | top_46_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1576_out | top_46_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? down_36_write_out : '0;
  assign top_46_read_write_en = (!(par_done_reg780_out | top_46_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg928_out | top_46_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1073_out | top_46_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1210_out | top_46_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1333_out | top_46_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1436_out | top_46_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1516_out | top_46_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1576_out | top_46_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign pe_46_top = (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? top_46_read_out : '0;
  assign pe_46_left = (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? left_46_read_out : '0;
  assign pe_46_go = (!pe_46_done & (!(par_done_reg884_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1030_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1169_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1296_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1405_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1492_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1558_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1606_out | right_46_write_done & down_46_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign down_45_write_in = (pe_45_done & (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_45_down : '0;
  assign down_45_write_write_en = (pe_45_done & (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign right_45_write_in = (pe_45_done & (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_45_right : '0;
  assign right_45_write_write_en = (pe_45_done & (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign left_45_read_in = (!(par_done_reg679_out | left_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg827_out | left_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg975_out | left_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1118_out | left_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1251_out | left_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1368_out | left_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1463_out | left_45_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1536_out | left_45_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? right_44_write_out : '0;
  assign left_45_read_write_en = (!(par_done_reg679_out | left_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg827_out | left_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg975_out | left_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1118_out | left_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1251_out | left_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1368_out | left_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1463_out | left_45_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1536_out | left_45_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign top_45_read_in = (!(par_done_reg633_out | top_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg779_out | top_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg927_out | top_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1072_out | top_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1209_out | top_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1332_out | top_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1435_out | top_45_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1515_out | top_45_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? down_35_write_out : '0;
  assign top_45_read_write_en = (!(par_done_reg633_out | top_45_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg779_out | top_45_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg927_out | top_45_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1072_out | top_45_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1209_out | top_45_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1332_out | top_45_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1435_out | top_45_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1515_out | top_45_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign pe_45_top = (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? top_45_read_out : '0;
  assign pe_45_left = (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? left_45_read_out : '0;
  assign pe_45_go = (!pe_45_done & (!(par_done_reg735_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg883_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1029_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1168_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1295_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1404_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1491_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1557_out | right_45_write_done & down_45_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign down_44_write_in = (pe_44_done & (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_44_down : '0;
  assign down_44_write_write_en = (pe_44_done & (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_44_write_in = (pe_44_done & (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_44_right : '0;
  assign right_44_write_write_en = (pe_44_done & (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_44_read_in = (!(par_done_reg536_out | left_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg678_out | left_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg826_out | left_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg974_out | left_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1117_out | left_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1250_out | left_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1367_out | left_44_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1462_out | left_44_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_43_write_out : '0;
  assign left_44_read_write_en = (!(par_done_reg536_out | left_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg678_out | left_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg826_out | left_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg974_out | left_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1117_out | left_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1250_out | left_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1367_out | left_44_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1462_out | left_44_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_44_read_in = (!(par_done_reg494_out | top_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg632_out | top_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg778_out | top_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg926_out | top_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1071_out | top_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1208_out | top_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1331_out | top_44_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1434_out | top_44_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_34_write_out : '0;
  assign top_44_read_write_en = (!(par_done_reg494_out | top_44_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg632_out | top_44_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg778_out | top_44_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg926_out | top_44_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1071_out | top_44_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1208_out | top_44_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1331_out | top_44_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1434_out | top_44_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_44_top = (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_44_read_out : '0;
  assign pe_44_left = (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_44_read_out : '0;
  assign pe_44_go = (!pe_44_done & (!(par_done_reg590_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg734_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg882_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1028_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1167_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1294_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1403_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1490_out | right_44_write_done & down_44_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign down_43_write_in = (pe_43_done & (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_43_down : '0;
  assign down_43_write_write_en = (pe_43_done & (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_43_write_in = (pe_43_done & (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_43_right : '0;
  assign right_43_write_write_en = (pe_43_done & (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_43_read_in = (!(par_done_reg405_out | left_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg535_out | left_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg677_out | left_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg825_out | left_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg973_out | left_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1116_out | left_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1249_out | left_43_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1366_out | left_43_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_42_write_out : '0;
  assign left_43_read_write_en = (!(par_done_reg405_out | left_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg535_out | left_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg677_out | left_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg825_out | left_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg973_out | left_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1116_out | left_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1249_out | left_43_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1366_out | left_43_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_43_read_in = (!(par_done_reg369_out | top_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg493_out | top_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg631_out | top_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg777_out | top_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg925_out | top_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1070_out | top_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1207_out | top_43_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1330_out | top_43_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_33_write_out : '0;
  assign top_43_read_write_en = (!(par_done_reg369_out | top_43_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg493_out | top_43_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg631_out | top_43_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg777_out | top_43_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg925_out | top_43_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1070_out | top_43_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1207_out | top_43_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1330_out | top_43_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_43_top = (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_43_read_out : '0;
  assign pe_43_left = (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_43_read_out : '0;
  assign pe_43_go = (!pe_43_done & (!(par_done_reg455_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg589_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg733_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg881_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1027_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1166_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1293_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1402_out | right_43_write_done & down_43_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_42_write_in = (pe_42_done & (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_42_down : '0;
  assign down_42_write_write_en = (pe_42_done & (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_42_write_in = (pe_42_done & (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_42_right : '0;
  assign right_42_write_write_en = (pe_42_done & (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_42_read_in = (!(par_done_reg292_out | left_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg404_out | left_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg534_out | left_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg676_out | left_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg824_out | left_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg972_out | left_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1115_out | left_42_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1248_out | left_42_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_41_write_out : '0;
  assign left_42_read_write_en = (!(par_done_reg292_out | left_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg404_out | left_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg534_out | left_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg676_out | left_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg824_out | left_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg972_out | left_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1115_out | left_42_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1248_out | left_42_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_42_read_in = (!(par_done_reg264_out | top_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg368_out | top_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg492_out | top_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg630_out | top_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg776_out | top_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg924_out | top_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1069_out | top_42_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1206_out | top_42_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_32_write_out : '0;
  assign top_42_read_write_en = (!(par_done_reg264_out | top_42_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg368_out | top_42_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg492_out | top_42_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg630_out | top_42_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg776_out | top_42_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg924_out | top_42_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1069_out | top_42_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1206_out | top_42_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_42_top = (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_42_read_out : '0;
  assign pe_42_left = (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_42_read_out : '0;
  assign pe_42_go = (!pe_42_done & (!(par_done_reg336_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg454_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg588_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg732_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg880_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1026_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1165_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1292_out | right_42_write_done & down_42_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_41_write_in = (pe_41_done & (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_41_down : '0;
  assign down_41_write_write_en = (pe_41_done & (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_41_write_in = (pe_41_done & (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_41_right : '0;
  assign right_41_write_write_en = (pe_41_done & (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_41_read_in = (!(par_done_reg203_out | left_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg291_out | left_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg403_out | left_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg533_out | left_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg675_out | left_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg823_out | left_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg971_out | left_41_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1114_out | left_41_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_40_write_out : '0;
  assign left_41_read_write_en = (!(par_done_reg203_out | left_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg291_out | left_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg403_out | left_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg533_out | left_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg675_out | left_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg823_out | left_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg971_out | left_41_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1114_out | left_41_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_41_read_in = (!(par_done_reg182_out | top_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg263_out | top_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg367_out | top_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg491_out | top_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg629_out | top_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg775_out | top_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg923_out | top_41_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1068_out | top_41_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_31_write_out : '0;
  assign top_41_read_write_en = (!(par_done_reg182_out | top_41_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg263_out | top_41_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg367_out | top_41_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg491_out | top_41_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg629_out | top_41_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg775_out | top_41_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg923_out | top_41_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1068_out | top_41_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_41_top = (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_41_read_out : '0;
  assign pe_41_left = (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_41_read_out : '0;
  assign pe_41_go = (!pe_41_done & (!(par_done_reg238_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg335_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg453_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg587_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg731_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg879_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1025_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1164_out | right_41_write_done & down_41_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_40_write_in = (pe_40_done & (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_40_down : '0;
  assign down_40_write_write_en = (pe_40_done & (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_40_write_in = (pe_40_done & (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_40_right : '0;
  assign right_40_write_write_en = (pe_40_done & (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_40_read_in = (!(par_done_reg135_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg202_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg290_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg402_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg532_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg674_out | left_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg822_out | left_40_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg970_out | left_40_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? l4_read_data : '0;
  assign left_40_read_write_en = (!(par_done_reg135_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg202_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg290_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg402_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg532_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg674_out | left_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg822_out | left_40_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg970_out | left_40_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_40_read_in = (!(par_done_reg120_out | top_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg181_out | top_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg262_out | top_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg366_out | top_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg490_out | top_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg628_out | top_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg774_out | top_40_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg922_out | top_40_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_30_write_out : '0;
  assign top_40_read_write_en = (!(par_done_reg120_out | top_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg181_out | top_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg262_out | top_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg366_out | top_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg490_out | top_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg628_out | top_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg774_out | top_40_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg922_out | top_40_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_40_top = (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_40_read_out : '0;
  assign pe_40_left = (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_40_read_out : '0;
  assign pe_40_go = (!pe_40_done & (!(par_done_reg162_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg237_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg334_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg452_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg586_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg730_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg878_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1024_out | right_40_write_done & down_40_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_37_write_in = (pe_37_done & (!(par_done_reg877_out | down_37_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1023_out | down_37_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1163_out | down_37_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1291_out | down_37_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1401_out | down_37_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1489_out | down_37_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1556_out | down_37_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1605_out | down_37_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? pe_37_down : '0;
  assign down_37_write_write_en = (pe_37_done & (!(par_done_reg877_out | down_37_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1023_out | down_37_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1163_out | down_37_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1291_out | down_37_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1401_out | down_37_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1489_out | down_37_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1556_out | down_37_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1605_out | down_37_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign left_37_read_in = (!(par_done_reg821_out | left_37_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg969_out | left_37_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1113_out | left_37_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1247_out | left_37_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1365_out | left_37_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1461_out | left_37_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1535_out | left_37_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1590_out | left_37_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? right_36_write_out : '0;
  assign left_37_read_write_en = (!(par_done_reg821_out | left_37_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg969_out | left_37_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1113_out | left_37_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1247_out | left_37_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1365_out | left_37_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1461_out | left_37_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1535_out | left_37_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1590_out | left_37_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign top_37_read_in = (!(par_done_reg773_out | top_37_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg921_out | top_37_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1067_out | top_37_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1205_out | top_37_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1329_out | top_37_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1433_out | top_37_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1514_out | top_37_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1575_out | top_37_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? down_27_write_out : '0;
  assign top_37_read_write_en = (!(par_done_reg773_out | top_37_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg921_out | top_37_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1067_out | top_37_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1205_out | top_37_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1329_out | top_37_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1433_out | top_37_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1514_out | top_37_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go | !(par_done_reg1575_out | top_37_read_done) & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign pe_37_top = (!(par_done_reg877_out | down_37_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1023_out | down_37_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1163_out | down_37_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1291_out | down_37_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1401_out | down_37_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1489_out | down_37_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1556_out | down_37_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1605_out | down_37_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? top_37_read_out : '0;
  assign pe_37_left = (!(par_done_reg877_out | down_37_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1023_out | down_37_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1163_out | down_37_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1291_out | down_37_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1401_out | down_37_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1489_out | down_37_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1556_out | down_37_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1605_out | down_37_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go) ? left_37_read_out : '0;
  assign pe_37_go = (!pe_37_done & (!(par_done_reg877_out | down_37_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1023_out | down_37_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1163_out | down_37_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1291_out | down_37_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1401_out | down_37_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1489_out | down_37_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1556_out | down_37_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go | !(par_done_reg1605_out | down_37_write_done) & fsm0_out == 32'd37 & !par_reset37_out & go)) ? 1'd1 : '0;
  assign down_36_write_in = (pe_36_done & (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_36_down : '0;
  assign down_36_write_write_en = (pe_36_done & (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign right_36_write_in = (pe_36_done & (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_36_right : '0;
  assign right_36_write_write_en = (pe_36_done & (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign left_36_read_in = (!(par_done_reg673_out | left_36_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg820_out | left_36_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg968_out | left_36_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1112_out | left_36_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1246_out | left_36_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1364_out | left_36_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1460_out | left_36_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1534_out | left_36_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? right_35_write_out : '0;
  assign left_36_read_write_en = (!(par_done_reg673_out | left_36_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg820_out | left_36_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg968_out | left_36_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1112_out | left_36_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1246_out | left_36_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1364_out | left_36_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1460_out | left_36_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1534_out | left_36_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign top_36_read_in = (!(par_done_reg627_out | top_36_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg772_out | top_36_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg920_out | top_36_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1066_out | top_36_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1204_out | top_36_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1328_out | top_36_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1432_out | top_36_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1513_out | top_36_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? down_26_write_out : '0;
  assign top_36_read_write_en = (!(par_done_reg627_out | top_36_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg772_out | top_36_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg920_out | top_36_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1066_out | top_36_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1204_out | top_36_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1328_out | top_36_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1432_out | top_36_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1513_out | top_36_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign pe_36_top = (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? top_36_read_out : '0;
  assign pe_36_left = (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? left_36_read_out : '0;
  assign pe_36_go = (!pe_36_done & (!(par_done_reg729_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg876_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1022_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1162_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1290_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1400_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1488_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1555_out | right_36_write_done & down_36_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign down_35_write_in = (pe_35_done & (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_35_down : '0;
  assign down_35_write_write_en = (pe_35_done & (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_35_write_in = (pe_35_done & (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_35_right : '0;
  assign right_35_write_write_en = (pe_35_done & (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_35_read_in = (!(par_done_reg531_out | left_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg672_out | left_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg819_out | left_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg967_out | left_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1111_out | left_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1245_out | left_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1363_out | left_35_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1459_out | left_35_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_34_write_out : '0;
  assign left_35_read_write_en = (!(par_done_reg531_out | left_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg672_out | left_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg819_out | left_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg967_out | left_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1111_out | left_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1245_out | left_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1363_out | left_35_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1459_out | left_35_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_35_read_in = (!(par_done_reg489_out | top_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg626_out | top_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg771_out | top_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg919_out | top_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1065_out | top_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1203_out | top_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1327_out | top_35_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1431_out | top_35_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_25_write_out : '0;
  assign top_35_read_write_en = (!(par_done_reg489_out | top_35_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg626_out | top_35_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg771_out | top_35_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg919_out | top_35_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1065_out | top_35_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1203_out | top_35_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1327_out | top_35_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1431_out | top_35_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_35_top = (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_35_read_out : '0;
  assign pe_35_left = (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_35_read_out : '0;
  assign pe_35_go = (!pe_35_done & (!(par_done_reg585_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg728_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg875_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1021_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1161_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1289_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1399_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1487_out | right_35_write_done & down_35_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign down_34_write_in = (pe_34_done & (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_34_down : '0;
  assign down_34_write_write_en = (pe_34_done & (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_34_write_in = (pe_34_done & (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_34_right : '0;
  assign right_34_write_write_en = (pe_34_done & (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_34_read_in = (!(par_done_reg401_out | left_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg530_out | left_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg671_out | left_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg818_out | left_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg966_out | left_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1110_out | left_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1244_out | left_34_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1362_out | left_34_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_33_write_out : '0;
  assign left_34_read_write_en = (!(par_done_reg401_out | left_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg530_out | left_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg671_out | left_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg818_out | left_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg966_out | left_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1110_out | left_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1244_out | left_34_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1362_out | left_34_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_34_read_in = (!(par_done_reg365_out | top_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg488_out | top_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg625_out | top_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg770_out | top_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg918_out | top_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1064_out | top_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1202_out | top_34_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1326_out | top_34_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_24_write_out : '0;
  assign top_34_read_write_en = (!(par_done_reg365_out | top_34_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg488_out | top_34_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg625_out | top_34_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg770_out | top_34_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg918_out | top_34_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1064_out | top_34_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1202_out | top_34_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1326_out | top_34_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_34_top = (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_34_read_out : '0;
  assign pe_34_left = (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_34_read_out : '0;
  assign pe_34_go = (!pe_34_done & (!(par_done_reg451_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg584_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg727_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg874_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1020_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1160_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1288_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1398_out | right_34_write_done & down_34_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_33_write_in = (pe_33_done & (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_33_down : '0;
  assign down_33_write_write_en = (pe_33_done & (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_33_write_in = (pe_33_done & (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_33_right : '0;
  assign right_33_write_write_en = (pe_33_done & (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_33_read_in = (!(par_done_reg289_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg400_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg529_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg670_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg817_out | left_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg965_out | left_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1109_out | left_33_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1243_out | left_33_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_32_write_out : '0;
  assign left_33_read_write_en = (!(par_done_reg289_out | left_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg400_out | left_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg529_out | left_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg670_out | left_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg817_out | left_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg965_out | left_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1109_out | left_33_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1243_out | left_33_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_33_read_in = (!(par_done_reg261_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg364_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg487_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg624_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg769_out | top_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg917_out | top_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1063_out | top_33_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1201_out | top_33_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_23_write_out : '0;
  assign top_33_read_write_en = (!(par_done_reg261_out | top_33_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg364_out | top_33_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg487_out | top_33_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg624_out | top_33_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg769_out | top_33_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg917_out | top_33_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1063_out | top_33_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1201_out | top_33_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_33_top = (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_33_read_out : '0;
  assign pe_33_left = (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_33_read_out : '0;
  assign pe_33_go = (!pe_33_done & (!(par_done_reg333_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg450_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg583_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg726_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg873_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1019_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1159_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1287_out | right_33_write_done & down_33_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_32_write_in = (pe_32_done & (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_32_down : '0;
  assign down_32_write_write_en = (pe_32_done & (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_32_write_in = (pe_32_done & (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_32_right : '0;
  assign right_32_write_write_en = (pe_32_done & (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_32_read_in = (!(par_done_reg201_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg288_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg399_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg528_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg669_out | left_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg816_out | left_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg964_out | left_32_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1108_out | left_32_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_31_write_out : '0;
  assign left_32_read_write_en = (!(par_done_reg201_out | left_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg288_out | left_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg399_out | left_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg528_out | left_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg669_out | left_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg816_out | left_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg964_out | left_32_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1108_out | left_32_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_32_read_in = (!(par_done_reg180_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg260_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg363_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg486_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg623_out | top_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg768_out | top_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg916_out | top_32_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1062_out | top_32_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_22_write_out : '0;
  assign top_32_read_write_en = (!(par_done_reg180_out | top_32_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg260_out | top_32_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg363_out | top_32_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg486_out | top_32_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg623_out | top_32_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg768_out | top_32_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg916_out | top_32_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1062_out | top_32_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_32_top = (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_32_read_out : '0;
  assign pe_32_left = (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_32_read_out : '0;
  assign pe_32_go = (!pe_32_done & (!(par_done_reg236_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg332_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg449_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg582_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg725_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg872_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1018_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1158_out | right_32_write_done & down_32_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_31_write_in = (pe_31_done & (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_31_down : '0;
  assign down_31_write_write_en = (pe_31_done & (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_31_write_in = (pe_31_done & (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_31_right : '0;
  assign right_31_write_write_en = (pe_31_done & (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_31_read_in = (!(par_done_reg134_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg200_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg287_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg398_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg527_out | left_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg668_out | left_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg815_out | left_31_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg963_out | left_31_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_30_write_out : '0;
  assign left_31_read_write_en = (!(par_done_reg134_out | left_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg200_out | left_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg287_out | left_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg398_out | left_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg527_out | left_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg668_out | left_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg815_out | left_31_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg963_out | left_31_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_31_read_in = (!(par_done_reg119_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg179_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg259_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg362_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg485_out | top_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg622_out | top_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg767_out | top_31_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg915_out | top_31_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_21_write_out : '0;
  assign top_31_read_write_en = (!(par_done_reg119_out | top_31_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg179_out | top_31_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg259_out | top_31_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg362_out | top_31_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg485_out | top_31_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg622_out | top_31_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg767_out | top_31_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg915_out | top_31_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_31_top = (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_31_read_out : '0;
  assign pe_31_left = (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_31_read_out : '0;
  assign pe_31_go = (!pe_31_done & (!(par_done_reg161_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg235_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg331_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg448_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg581_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg724_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg871_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1017_out | right_31_write_done & down_31_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_30_write_in = (pe_30_done & (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_30_down : '0;
  assign down_30_write_write_en = (pe_30_done & (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_30_write_in = (pe_30_done & (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_30_right : '0;
  assign right_30_write_write_en = (pe_30_done & (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_30_read_in = (!(par_done_reg85_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg133_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg199_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg286_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg397_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg526_out | left_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg667_out | left_30_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg814_out | left_30_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? l3_read_data : '0;
  assign left_30_read_write_en = (!(par_done_reg85_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg133_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg199_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg286_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg397_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg526_out | left_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg667_out | left_30_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg814_out | left_30_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_30_read_in = (!(par_done_reg75_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg118_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg178_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg258_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg361_out | top_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg484_out | top_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg621_out | top_30_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg766_out | top_30_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_20_write_out : '0;
  assign top_30_read_write_en = (!(par_done_reg75_out | top_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg118_out | top_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg178_out | top_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg258_out | top_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg361_out | top_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg484_out | top_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg621_out | top_30_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg766_out | top_30_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_30_top = (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_30_read_out : '0;
  assign pe_30_left = (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_30_read_out : '0;
  assign pe_30_go = (!pe_30_done & (!(par_done_reg105_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg160_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg234_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg330_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg447_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg580_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg723_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg870_out | right_30_write_done & down_30_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_27_write_in = (pe_27_done & (!(par_done_reg722_out | down_27_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg869_out | down_27_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1016_out | down_27_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1157_out | down_27_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1286_out | down_27_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1397_out | down_27_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1486_out | down_27_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1554_out | down_27_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? pe_27_down : '0;
  assign down_27_write_write_en = (pe_27_done & (!(par_done_reg722_out | down_27_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg869_out | down_27_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1016_out | down_27_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1157_out | down_27_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1286_out | down_27_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1397_out | down_27_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1486_out | down_27_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1554_out | down_27_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign left_27_read_in = (!(par_done_reg666_out | left_27_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg813_out | left_27_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg962_out | left_27_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1107_out | left_27_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1242_out | left_27_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1361_out | left_27_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1458_out | left_27_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1533_out | left_27_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? right_26_write_out : '0;
  assign left_27_read_write_en = (!(par_done_reg666_out | left_27_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg813_out | left_27_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg962_out | left_27_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1107_out | left_27_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1242_out | left_27_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1361_out | left_27_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1458_out | left_27_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1533_out | left_27_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign top_27_read_in = (!(par_done_reg620_out | top_27_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg765_out | top_27_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg914_out | top_27_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1061_out | top_27_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1200_out | top_27_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1325_out | top_27_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1430_out | top_27_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1512_out | top_27_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? down_17_write_out : '0;
  assign top_27_read_write_en = (!(par_done_reg620_out | top_27_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg765_out | top_27_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg914_out | top_27_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1061_out | top_27_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1200_out | top_27_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1325_out | top_27_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1430_out | top_27_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go | !(par_done_reg1512_out | top_27_read_done) & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign pe_27_top = (!(par_done_reg722_out | down_27_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg869_out | down_27_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1016_out | down_27_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1157_out | down_27_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1286_out | down_27_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1397_out | down_27_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1486_out | down_27_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1554_out | down_27_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? top_27_read_out : '0;
  assign pe_27_left = (!(par_done_reg722_out | down_27_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg869_out | down_27_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1016_out | down_27_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1157_out | down_27_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1286_out | down_27_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1397_out | down_27_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1486_out | down_27_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1554_out | down_27_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go) ? left_27_read_out : '0;
  assign pe_27_go = (!pe_27_done & (!(par_done_reg722_out | down_27_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg869_out | down_27_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1016_out | down_27_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1157_out | down_27_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1286_out | down_27_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1397_out | down_27_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1486_out | down_27_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go | !(par_done_reg1554_out | down_27_write_done) & fsm0_out == 32'd35 & !par_reset35_out & go)) ? 1'd1 : '0;
  assign down_26_write_in = (pe_26_done & (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_26_down : '0;
  assign down_26_write_write_en = (pe_26_done & (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign right_26_write_in = (pe_26_done & (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_26_right : '0;
  assign right_26_write_write_en = (pe_26_done & (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_26_read_in = (!(par_done_reg525_out | left_26_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg665_out | left_26_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg812_out | left_26_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg961_out | left_26_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1106_out | left_26_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1241_out | left_26_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1360_out | left_26_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1457_out | left_26_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_25_write_out : '0;
  assign left_26_read_write_en = (!(par_done_reg525_out | left_26_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg665_out | left_26_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg812_out | left_26_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg961_out | left_26_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1106_out | left_26_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1241_out | left_26_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1360_out | left_26_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1457_out | left_26_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_26_read_in = (!(par_done_reg483_out | top_26_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg619_out | top_26_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg764_out | top_26_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg913_out | top_26_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1060_out | top_26_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1199_out | top_26_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1324_out | top_26_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1429_out | top_26_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_16_write_out : '0;
  assign top_26_read_write_en = (!(par_done_reg483_out | top_26_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg619_out | top_26_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg764_out | top_26_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg913_out | top_26_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1060_out | top_26_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1199_out | top_26_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1324_out | top_26_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1429_out | top_26_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_26_top = (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_26_read_out : '0;
  assign pe_26_left = (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_26_read_out : '0;
  assign pe_26_go = (!pe_26_done & (!(par_done_reg579_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg721_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg868_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1015_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1156_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1285_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1396_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1485_out | right_26_write_done & down_26_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign down_25_write_in = (pe_25_done & (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_25_down : '0;
  assign down_25_write_write_en = (pe_25_done & (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_25_write_in = (pe_25_done & (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_25_right : '0;
  assign right_25_write_write_en = (pe_25_done & (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_25_read_in = (!(par_done_reg396_out | left_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg524_out | left_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg664_out | left_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg811_out | left_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg960_out | left_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1105_out | left_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1240_out | left_25_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1359_out | left_25_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_24_write_out : '0;
  assign left_25_read_write_en = (!(par_done_reg396_out | left_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg524_out | left_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg664_out | left_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg811_out | left_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg960_out | left_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1105_out | left_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1240_out | left_25_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1359_out | left_25_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_25_read_in = (!(par_done_reg360_out | top_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg482_out | top_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg618_out | top_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg763_out | top_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg912_out | top_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1059_out | top_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1198_out | top_25_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1323_out | top_25_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_15_write_out : '0;
  assign top_25_read_write_en = (!(par_done_reg360_out | top_25_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg482_out | top_25_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg618_out | top_25_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg763_out | top_25_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg912_out | top_25_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1059_out | top_25_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1198_out | top_25_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1323_out | top_25_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_25_top = (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_25_read_out : '0;
  assign pe_25_left = (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_25_read_out : '0;
  assign pe_25_go = (!pe_25_done & (!(par_done_reg446_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg578_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg720_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg867_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1014_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1155_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1284_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1395_out | right_25_write_done & down_25_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_24_write_in = (pe_24_done & (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_24_down : '0;
  assign down_24_write_write_en = (pe_24_done & (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_24_write_in = (pe_24_done & (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_24_right : '0;
  assign right_24_write_write_en = (pe_24_done & (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_24_read_in = (!(par_done_reg285_out | left_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg395_out | left_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg523_out | left_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg663_out | left_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg810_out | left_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg959_out | left_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1104_out | left_24_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1239_out | left_24_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_23_write_out : '0;
  assign left_24_read_write_en = (!(par_done_reg285_out | left_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg395_out | left_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg523_out | left_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg663_out | left_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg810_out | left_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg959_out | left_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1104_out | left_24_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1239_out | left_24_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_24_read_in = (!(par_done_reg257_out | top_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg359_out | top_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg481_out | top_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg617_out | top_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg762_out | top_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg911_out | top_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1058_out | top_24_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1197_out | top_24_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_14_write_out : '0;
  assign top_24_read_write_en = (!(par_done_reg257_out | top_24_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg359_out | top_24_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg481_out | top_24_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg617_out | top_24_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg762_out | top_24_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg911_out | top_24_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1058_out | top_24_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1197_out | top_24_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_24_top = (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_24_read_out : '0;
  assign pe_24_left = (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_24_read_out : '0;
  assign pe_24_go = (!pe_24_done & (!(par_done_reg329_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg445_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg577_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg719_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg866_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1013_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1154_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1283_out | right_24_write_done & down_24_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_23_write_in = (pe_23_done & (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_23_down : '0;
  assign down_23_write_write_en = (pe_23_done & (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_23_write_in = (pe_23_done & (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_23_right : '0;
  assign right_23_write_write_en = (pe_23_done & (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_23_read_in = (!(par_done_reg198_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg284_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg394_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg522_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg662_out | left_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg809_out | left_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg958_out | left_23_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1103_out | left_23_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_22_write_out : '0;
  assign left_23_read_write_en = (!(par_done_reg198_out | left_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg284_out | left_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg394_out | left_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg522_out | left_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg662_out | left_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg809_out | left_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg958_out | left_23_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1103_out | left_23_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_23_read_in = (!(par_done_reg177_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg256_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg358_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg480_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg616_out | top_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg761_out | top_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg910_out | top_23_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1057_out | top_23_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_13_write_out : '0;
  assign top_23_read_write_en = (!(par_done_reg177_out | top_23_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg256_out | top_23_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg358_out | top_23_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg480_out | top_23_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg616_out | top_23_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg761_out | top_23_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg910_out | top_23_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1057_out | top_23_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_23_top = (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_23_read_out : '0;
  assign pe_23_left = (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_23_read_out : '0;
  assign pe_23_go = (!pe_23_done & (!(par_done_reg233_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg328_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg444_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg576_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg718_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg865_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1012_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1153_out | right_23_write_done & down_23_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_22_write_in = (pe_22_done & (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_22_down : '0;
  assign down_22_write_write_en = (pe_22_done & (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_22_write_in = (pe_22_done & (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_22_right : '0;
  assign right_22_write_write_en = (pe_22_done & (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_22_read_in = (!(par_done_reg132_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg197_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg283_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg393_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg521_out | left_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg661_out | left_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg808_out | left_22_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg957_out | left_22_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_21_write_out : '0;
  assign left_22_read_write_en = (!(par_done_reg132_out | left_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg197_out | left_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg283_out | left_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg393_out | left_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg521_out | left_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg661_out | left_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg808_out | left_22_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg957_out | left_22_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_22_read_in = (!(par_done_reg117_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg176_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg255_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg357_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg479_out | top_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg615_out | top_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg760_out | top_22_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg909_out | top_22_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_12_write_out : '0;
  assign top_22_read_write_en = (!(par_done_reg117_out | top_22_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg176_out | top_22_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg255_out | top_22_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg357_out | top_22_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg479_out | top_22_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg615_out | top_22_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg760_out | top_22_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg909_out | top_22_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_22_top = (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_22_read_out : '0;
  assign pe_22_left = (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_22_read_out : '0;
  assign pe_22_go = (!pe_22_done & (!(par_done_reg159_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg232_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg327_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg443_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg575_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg717_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg864_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1011_out | right_22_write_done & down_22_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_21_write_in = (pe_21_done & (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_21_down : '0;
  assign down_21_write_write_en = (pe_21_done & (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_21_write_in = (pe_21_done & (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_21_right : '0;
  assign right_21_write_write_en = (pe_21_done & (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_21_read_in = (!(par_done_reg84_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg131_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg196_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg282_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg392_out | left_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg520_out | left_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg660_out | left_21_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg807_out | left_21_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_20_write_out : '0;
  assign left_21_read_write_en = (!(par_done_reg84_out | left_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg131_out | left_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg196_out | left_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg282_out | left_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg392_out | left_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg520_out | left_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg660_out | left_21_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg807_out | left_21_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_21_read_in = (!(par_done_reg74_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg254_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg356_out | top_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg478_out | top_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg614_out | top_21_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg759_out | top_21_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_11_write_out : '0;
  assign top_21_read_write_en = (!(par_done_reg74_out | top_21_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg116_out | top_21_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg175_out | top_21_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg254_out | top_21_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg356_out | top_21_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg478_out | top_21_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg614_out | top_21_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg759_out | top_21_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_21_top = (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_21_read_out : '0;
  assign pe_21_left = (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_21_read_out : '0;
  assign pe_21_go = (!pe_21_done & (!(par_done_reg104_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg158_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg231_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg326_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg442_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg574_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg716_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg863_out | right_21_write_done & down_21_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_20_write_in = (pe_20_done & (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_20_down : '0;
  assign down_20_write_write_en = (pe_20_done & (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_20_write_in = (pe_20_done & (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_20_right : '0;
  assign right_20_write_write_en = (pe_20_done & (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_20_read_in = (!(par_done_reg51_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg83_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg130_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg195_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg281_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg391_out | left_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg519_out | left_20_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg659_out | left_20_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? l2_read_data : '0;
  assign left_20_read_write_en = (!(par_done_reg51_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg83_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg130_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg195_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg281_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg391_out | left_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg519_out | left_20_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg659_out | left_20_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_20_read_in = (!(par_done_reg45_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg73_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg115_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg174_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg253_out | top_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg355_out | top_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg477_out | top_20_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg613_out | top_20_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_10_write_out : '0;
  assign top_20_read_write_en = (!(par_done_reg45_out | top_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg73_out | top_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg115_out | top_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg174_out | top_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg253_out | top_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg355_out | top_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg477_out | top_20_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg613_out | top_20_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_20_top = (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_20_read_out : '0;
  assign pe_20_left = (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_20_read_out : '0;
  assign pe_20_go = (!pe_20_done & (!(par_done_reg65_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg103_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg157_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg230_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg325_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg441_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg573_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg715_out | right_20_write_done & down_20_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_17_write_in = (pe_17_done & (!(par_done_reg572_out | down_17_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg714_out | down_17_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg862_out | down_17_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1010_out | down_17_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1152_out | down_17_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1282_out | down_17_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1394_out | down_17_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1484_out | down_17_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? pe_17_down : '0;
  assign down_17_write_write_en = (pe_17_done & (!(par_done_reg572_out | down_17_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg714_out | down_17_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg862_out | down_17_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1010_out | down_17_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1152_out | down_17_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1282_out | down_17_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1394_out | down_17_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1484_out | down_17_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign left_17_read_in = (!(par_done_reg518_out | left_17_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg658_out | left_17_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg806_out | left_17_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg956_out | left_17_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1102_out | left_17_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1238_out | left_17_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1358_out | left_17_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1456_out | left_17_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? right_16_write_out : '0;
  assign left_17_read_write_en = (!(par_done_reg518_out | left_17_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg658_out | left_17_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg806_out | left_17_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg956_out | left_17_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1102_out | left_17_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1238_out | left_17_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1358_out | left_17_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1456_out | left_17_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign top_17_read_in = (!(par_done_reg476_out | top_17_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg612_out | top_17_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg758_out | top_17_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg908_out | top_17_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1056_out | top_17_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1196_out | top_17_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1322_out | top_17_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1428_out | top_17_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? down_07_write_out : '0;
  assign top_17_read_write_en = (!(par_done_reg476_out | top_17_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg612_out | top_17_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg758_out | top_17_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg908_out | top_17_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1056_out | top_17_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1196_out | top_17_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1322_out | top_17_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go | !(par_done_reg1428_out | top_17_read_done) & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign pe_17_top = (!(par_done_reg572_out | down_17_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg714_out | down_17_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg862_out | down_17_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1010_out | down_17_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1152_out | down_17_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1282_out | down_17_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1394_out | down_17_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1484_out | down_17_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? top_17_read_out : '0;
  assign pe_17_left = (!(par_done_reg572_out | down_17_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg714_out | down_17_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg862_out | down_17_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1010_out | down_17_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1152_out | down_17_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1282_out | down_17_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1394_out | down_17_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1484_out | down_17_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go) ? left_17_read_out : '0;
  assign pe_17_go = (!pe_17_done & (!(par_done_reg572_out | down_17_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg714_out | down_17_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg862_out | down_17_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1010_out | down_17_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1152_out | down_17_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1282_out | down_17_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1394_out | down_17_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go | !(par_done_reg1484_out | down_17_write_done) & fsm0_out == 32'd33 & !par_reset33_out & go)) ? 1'd1 : '0;
  assign down_16_write_in = (pe_16_done & (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_16_down : '0;
  assign down_16_write_write_en = (pe_16_done & (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign right_16_write_in = (pe_16_done & (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_16_right : '0;
  assign right_16_write_write_en = (pe_16_done & (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_16_read_in = (!(par_done_reg390_out | left_16_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg517_out | left_16_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg657_out | left_16_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg805_out | left_16_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg955_out | left_16_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1101_out | left_16_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1237_out | left_16_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1357_out | left_16_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_15_write_out : '0;
  assign left_16_read_write_en = (!(par_done_reg390_out | left_16_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg517_out | left_16_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg657_out | left_16_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg805_out | left_16_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg955_out | left_16_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1101_out | left_16_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1237_out | left_16_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1357_out | left_16_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_16_read_in = (!(par_done_reg354_out | top_16_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg475_out | top_16_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg611_out | top_16_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg757_out | top_16_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg907_out | top_16_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1055_out | top_16_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1195_out | top_16_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1321_out | top_16_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? down_06_write_out : '0;
  assign top_16_read_write_en = (!(par_done_reg354_out | top_16_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg475_out | top_16_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg611_out | top_16_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg757_out | top_16_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg907_out | top_16_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1055_out | top_16_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1195_out | top_16_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1321_out | top_16_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_16_top = (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_16_read_out : '0;
  assign pe_16_left = (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_16_read_out : '0;
  assign pe_16_go = (!pe_16_done & (!(par_done_reg440_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg571_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg713_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg861_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1009_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1151_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1281_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1393_out | right_16_write_done & down_16_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_15_write_in = (pe_15_done & (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_15_down : '0;
  assign down_15_write_write_en = (pe_15_done & (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_15_write_in = (pe_15_done & (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_15_right : '0;
  assign right_15_write_write_en = (pe_15_done & (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_15_read_in = (!(par_done_reg280_out | left_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg389_out | left_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg516_out | left_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg656_out | left_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg804_out | left_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg954_out | left_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1100_out | left_15_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1236_out | left_15_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_14_write_out : '0;
  assign left_15_read_write_en = (!(par_done_reg280_out | left_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg389_out | left_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg516_out | left_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg656_out | left_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg804_out | left_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg954_out | left_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1100_out | left_15_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1236_out | left_15_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_15_read_in = (!(par_done_reg252_out | top_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg353_out | top_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg474_out | top_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg610_out | top_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg756_out | top_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg906_out | top_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1054_out | top_15_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1194_out | top_15_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? down_05_write_out : '0;
  assign top_15_read_write_en = (!(par_done_reg252_out | top_15_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg353_out | top_15_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg474_out | top_15_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg610_out | top_15_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg756_out | top_15_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg906_out | top_15_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1054_out | top_15_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1194_out | top_15_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_15_top = (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_15_read_out : '0;
  assign pe_15_left = (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_15_read_out : '0;
  assign pe_15_go = (!pe_15_done & (!(par_done_reg324_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg439_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg570_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg712_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg860_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1008_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1150_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1280_out | right_15_write_done & down_15_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_14_write_in = (pe_14_done & (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_14_down : '0;
  assign down_14_write_write_en = (pe_14_done & (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_14_write_in = (pe_14_done & (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_14_right : '0;
  assign right_14_write_write_en = (pe_14_done & (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_14_read_in = (!(par_done_reg194_out | left_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg279_out | left_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg388_out | left_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg515_out | left_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg655_out | left_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg803_out | left_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg953_out | left_14_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1099_out | left_14_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_13_write_out : '0;
  assign left_14_read_write_en = (!(par_done_reg194_out | left_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg279_out | left_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg388_out | left_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg515_out | left_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg655_out | left_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg803_out | left_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg953_out | left_14_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1099_out | left_14_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_14_read_in = (!(par_done_reg173_out | top_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg251_out | top_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg352_out | top_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg473_out | top_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg609_out | top_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg755_out | top_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg905_out | top_14_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1053_out | top_14_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? down_04_write_out : '0;
  assign top_14_read_write_en = (!(par_done_reg173_out | top_14_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg251_out | top_14_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg352_out | top_14_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg473_out | top_14_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg609_out | top_14_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg755_out | top_14_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg905_out | top_14_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1053_out | top_14_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_14_top = (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_14_read_out : '0;
  assign pe_14_left = (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_14_read_out : '0;
  assign pe_14_go = (!pe_14_done & (!(par_done_reg229_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg323_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg438_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg569_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg711_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg859_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1007_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1149_out | right_14_write_done & down_14_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_13_write_in = (pe_13_done & (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_13_down : '0;
  assign down_13_write_write_en = (pe_13_done & (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_13_write_in = (pe_13_done & (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_13_right : '0;
  assign right_13_write_write_en = (pe_13_done & (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_13_read_in = (!(par_done_reg129_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg193_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg278_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg387_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg514_out | left_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg654_out | left_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg802_out | left_13_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg952_out | left_13_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_12_write_out : '0;
  assign left_13_read_write_en = (!(par_done_reg129_out | left_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg193_out | left_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg278_out | left_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg387_out | left_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg514_out | left_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg654_out | left_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg802_out | left_13_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg952_out | left_13_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_13_read_in = (!(par_done_reg114_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg172_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg250_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg351_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg472_out | top_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg608_out | top_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg754_out | top_13_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg904_out | top_13_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? down_03_write_out : '0;
  assign top_13_read_write_en = (!(par_done_reg114_out | top_13_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg172_out | top_13_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg250_out | top_13_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg351_out | top_13_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg472_out | top_13_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg608_out | top_13_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg754_out | top_13_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg904_out | top_13_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_13_top = (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_13_read_out : '0;
  assign pe_13_left = (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_13_read_out : '0;
  assign pe_13_go = (!pe_13_done & (!(par_done_reg156_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg228_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg322_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg437_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg568_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg710_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg858_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1006_out | right_13_write_done & down_13_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_12_write_in = (pe_12_done & (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_12_down : '0;
  assign down_12_write_write_en = (pe_12_done & (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_12_write_in = (pe_12_done & (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_12_right : '0;
  assign right_12_write_write_en = (pe_12_done & (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_12_read_in = (!(par_done_reg82_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg128_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg192_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg277_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg386_out | left_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg513_out | left_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg653_out | left_12_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg801_out | left_12_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_11_write_out : '0;
  assign left_12_read_write_en = (!(par_done_reg82_out | left_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg128_out | left_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg192_out | left_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg277_out | left_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg386_out | left_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg513_out | left_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg653_out | left_12_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg801_out | left_12_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_12_read_in = (!(par_done_reg72_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg113_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg171_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg249_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg350_out | top_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg471_out | top_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg607_out | top_12_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg753_out | top_12_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? down_02_write_out : '0;
  assign top_12_read_write_en = (!(par_done_reg72_out | top_12_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg113_out | top_12_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg171_out | top_12_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg249_out | top_12_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg350_out | top_12_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg471_out | top_12_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg607_out | top_12_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg753_out | top_12_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_12_top = (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_12_read_out : '0;
  assign pe_12_left = (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_12_read_out : '0;
  assign pe_12_go = (!pe_12_done & (!(par_done_reg102_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg155_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg227_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg321_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg436_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg567_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg709_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg857_out | right_12_write_done & down_12_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_11_write_in = (pe_11_done & (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_11_down : '0;
  assign down_11_write_write_en = (pe_11_done & (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_11_write_in = (pe_11_done & (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_11_right : '0;
  assign right_11_write_write_en = (pe_11_done & (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_11_read_in = (!(par_done_reg50_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg81_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg191_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg276_out | left_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg385_out | left_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg512_out | left_11_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg652_out | left_11_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_10_write_out : '0;
  assign left_11_read_write_en = (!(par_done_reg50_out | left_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg81_out | left_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg127_out | left_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg191_out | left_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg276_out | left_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg385_out | left_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg512_out | left_11_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg652_out | left_11_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_11_read_in = (!(par_done_reg44_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg71_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg112_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg170_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | top_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg349_out | top_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg470_out | top_11_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg606_out | top_11_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? down_01_write_out : '0;
  assign top_11_read_write_en = (!(par_done_reg44_out | top_11_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg71_out | top_11_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg112_out | top_11_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg170_out | top_11_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg248_out | top_11_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg349_out | top_11_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg470_out | top_11_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg606_out | top_11_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_11_top = (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_11_read_out : '0;
  assign pe_11_left = (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_11_read_out : '0;
  assign pe_11_go = (!pe_11_done & (!(par_done_reg64_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg101_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg154_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg226_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg320_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg435_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg566_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg708_out | right_11_write_done & down_11_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_10_write_in = (pe_10_done & (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_10_down : '0;
  assign down_10_write_write_en = (pe_10_done & (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_10_write_in = (pe_10_done & (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_10_right : '0;
  assign right_10_write_write_en = (pe_10_done & (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_10_read_in = (!(par_done_reg30_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg49_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg80_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg126_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg190_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg275_out | left_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg384_out | left_10_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg511_out | left_10_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? l1_read_data : '0;
  assign left_10_read_write_en = (!(par_done_reg30_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg49_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg80_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg126_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg190_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg275_out | left_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg384_out | left_10_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg511_out | left_10_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_10_read_in = (!(par_done_reg27_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg111_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg169_out | top_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg247_out | top_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg348_out | top_10_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg469_out | top_10_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? down_00_write_out : '0;
  assign top_10_read_write_en = (!(par_done_reg27_out | top_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg43_out | top_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg70_out | top_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg111_out | top_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg169_out | top_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg247_out | top_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg348_out | top_10_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg469_out | top_10_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_10_top = (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_10_read_out : '0;
  assign pe_10_left = (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_10_read_out : '0;
  assign pe_10_go = (!pe_10_done & (!(par_done_reg39_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg63_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg100_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg153_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg225_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg319_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg434_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg565_out | right_10_write_done & down_10_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_07_write_in = (pe_07_done & (!(par_done_reg433_out | down_07_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg564_out | down_07_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg707_out | down_07_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg856_out | down_07_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1005_out | down_07_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1148_out | down_07_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1279_out | down_07_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1392_out | down_07_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? pe_07_down : '0;
  assign down_07_write_write_en = (pe_07_done & (!(par_done_reg433_out | down_07_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg564_out | down_07_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg707_out | down_07_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg856_out | down_07_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1005_out | down_07_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1148_out | down_07_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1279_out | down_07_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1392_out | down_07_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign left_07_read_in = (!(par_done_reg383_out | left_07_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg510_out | left_07_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg651_out | left_07_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg800_out | left_07_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg951_out | left_07_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1098_out | left_07_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1235_out | left_07_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1356_out | left_07_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? right_06_write_out : '0;
  assign left_07_read_write_en = (!(par_done_reg383_out | left_07_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg510_out | left_07_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg651_out | left_07_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg800_out | left_07_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg951_out | left_07_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1098_out | left_07_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1235_out | left_07_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1356_out | left_07_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign top_07_read_in = (!(par_done_reg347_out | top_07_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg468_out | top_07_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg605_out | top_07_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg752_out | top_07_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg903_out | top_07_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1052_out | top_07_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1193_out | top_07_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1320_out | top_07_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? t7_read_data : '0;
  assign top_07_read_write_en = (!(par_done_reg347_out | top_07_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg468_out | top_07_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg605_out | top_07_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg752_out | top_07_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg903_out | top_07_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1052_out | top_07_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1193_out | top_07_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1320_out | top_07_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign pe_07_top = (!(par_done_reg433_out | down_07_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg564_out | down_07_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg707_out | down_07_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg856_out | down_07_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1005_out | down_07_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1148_out | down_07_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1279_out | down_07_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1392_out | down_07_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? top_07_read_out : '0;
  assign pe_07_left = (!(par_done_reg433_out | down_07_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg564_out | down_07_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg707_out | down_07_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg856_out | down_07_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1005_out | down_07_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1148_out | down_07_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1279_out | down_07_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1392_out | down_07_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go) ? left_07_read_out : '0;
  assign pe_07_go = (!pe_07_done & (!(par_done_reg433_out | down_07_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg564_out | down_07_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg707_out | down_07_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg856_out | down_07_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1005_out | down_07_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1148_out | down_07_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1279_out | down_07_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go | !(par_done_reg1392_out | down_07_write_done) & fsm0_out == 32'd31 & !par_reset31_out & go)) ? 1'd1 : '0;
  assign down_06_write_in = (pe_06_done & (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_06_down : '0;
  assign down_06_write_write_en = (pe_06_done & (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign right_06_write_in = (pe_06_done & (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? pe_06_right : '0;
  assign right_06_write_write_en = (pe_06_done & (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign left_06_read_in = (!(par_done_reg274_out | left_06_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg382_out | left_06_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg509_out | left_06_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg650_out | left_06_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg799_out | left_06_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg950_out | left_06_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1097_out | left_06_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1234_out | left_06_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? right_05_write_out : '0;
  assign left_06_read_write_en = (!(par_done_reg274_out | left_06_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg382_out | left_06_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg509_out | left_06_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg650_out | left_06_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg799_out | left_06_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg950_out | left_06_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1097_out | left_06_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1234_out | left_06_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign top_06_read_in = (!(par_done_reg246_out | top_06_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg346_out | top_06_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg467_out | top_06_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg604_out | top_06_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg751_out | top_06_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg902_out | top_06_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1051_out | top_06_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1192_out | top_06_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? t6_read_data : '0;
  assign top_06_read_write_en = (!(par_done_reg246_out | top_06_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg346_out | top_06_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg467_out | top_06_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg604_out | top_06_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg751_out | top_06_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg902_out | top_06_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1051_out | top_06_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1192_out | top_06_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign pe_06_top = (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? top_06_read_out : '0;
  assign pe_06_left = (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? left_06_read_out : '0;
  assign pe_06_go = (!pe_06_done & (!(par_done_reg318_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg432_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg563_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg706_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg855_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1004_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1147_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1278_out | right_06_write_done & down_06_write_done) & fsm0_out == 32'd29 & !par_reset29_out & go)) ? 1'd1 : '0;
  assign down_05_write_in = (pe_05_done & (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_05_down : '0;
  assign down_05_write_write_en = (pe_05_done & (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign right_05_write_in = (pe_05_done & (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? pe_05_right : '0;
  assign right_05_write_write_en = (pe_05_done & (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign left_05_read_in = (!(par_done_reg189_out | left_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg273_out | left_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg381_out | left_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg508_out | left_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg649_out | left_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg798_out | left_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg949_out | left_05_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1096_out | left_05_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? right_04_write_out : '0;
  assign left_05_read_write_en = (!(par_done_reg189_out | left_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg273_out | left_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg381_out | left_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg508_out | left_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg649_out | left_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg798_out | left_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg949_out | left_05_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1096_out | left_05_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign top_05_read_in = (!(par_done_reg168_out | top_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | top_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg345_out | top_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg466_out | top_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg603_out | top_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg750_out | top_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg901_out | top_05_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1050_out | top_05_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? t5_read_data : '0;
  assign top_05_read_write_en = (!(par_done_reg168_out | top_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | top_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg345_out | top_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg466_out | top_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg603_out | top_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg750_out | top_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg901_out | top_05_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1050_out | top_05_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign pe_05_top = (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? top_05_read_out : '0;
  assign pe_05_left = (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? left_05_read_out : '0;
  assign pe_05_go = (!pe_05_done & (!(par_done_reg224_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg317_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg431_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg562_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg705_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg854_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1003_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1146_out | right_05_write_done & down_05_write_done) & fsm0_out == 32'd27 & !par_reset27_out & go)) ? 1'd1 : '0;
  assign down_04_write_in = (pe_04_done & (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_04_down : '0;
  assign down_04_write_write_en = (pe_04_done & (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign right_04_write_in = (pe_04_done & (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? pe_04_right : '0;
  assign right_04_write_write_en = (pe_04_done & (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign left_04_read_in = (!(par_done_reg125_out | left_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg188_out | left_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg272_out | left_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg380_out | left_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg507_out | left_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg648_out | left_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg797_out | left_04_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg948_out | left_04_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? right_03_write_out : '0;
  assign left_04_read_write_en = (!(par_done_reg125_out | left_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg188_out | left_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg272_out | left_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg380_out | left_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg507_out | left_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg648_out | left_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg797_out | left_04_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg948_out | left_04_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign top_04_read_in = (!(par_done_reg110_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg344_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg465_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg602_out | top_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg749_out | top_04_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg900_out | top_04_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? t4_read_data : '0;
  assign top_04_read_write_en = (!(par_done_reg110_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg344_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg465_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg602_out | top_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg749_out | top_04_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg900_out | top_04_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign pe_04_top = (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? top_04_read_out : '0;
  assign pe_04_left = (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? left_04_read_out : '0;
  assign pe_04_go = (!pe_04_done & (!(par_done_reg152_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg223_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg316_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg430_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg561_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg704_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg853_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1002_out | right_04_write_done & down_04_write_done) & fsm0_out == 32'd25 & !par_reset25_out & go)) ? 1'd1 : '0;
  assign down_03_write_in = (pe_03_done & (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_03_down : '0;
  assign down_03_write_write_en = (pe_03_done & (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign right_03_write_in = (pe_03_done & (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? pe_03_right : '0;
  assign right_03_write_write_en = (pe_03_done & (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign left_03_read_in = (!(par_done_reg79_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg271_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg379_out | left_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg506_out | left_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg647_out | left_03_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg796_out | left_03_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? right_02_write_out : '0;
  assign left_03_read_write_en = (!(par_done_reg79_out | left_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg124_out | left_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg187_out | left_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg271_out | left_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg379_out | left_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg506_out | left_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg647_out | left_03_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg796_out | left_03_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign top_03_read_in = (!(par_done_reg69_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg243_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg343_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg464_out | top_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg601_out | top_03_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg748_out | top_03_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? t3_read_data : '0;
  assign top_03_read_write_en = (!(par_done_reg69_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg243_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg343_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg464_out | top_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg601_out | top_03_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg748_out | top_03_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign pe_03_top = (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? top_03_read_out : '0;
  assign pe_03_left = (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? left_03_read_out : '0;
  assign pe_03_go = (!pe_03_done & (!(par_done_reg99_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg151_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg222_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg315_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg429_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg560_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg703_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg852_out | right_03_write_done & down_03_write_done) & fsm0_out == 32'd23 & !par_reset23_out & go)) ? 1'd1 : '0;
  assign down_02_write_in = (pe_02_done & (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_02_down : '0;
  assign down_02_write_write_en = (pe_02_done & (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign right_02_write_in = (pe_02_done & (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? pe_02_right : '0;
  assign right_02_write_write_en = (pe_02_done & (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign left_02_read_in = (!(par_done_reg48_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg78_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg123_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg186_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg270_out | left_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg378_out | left_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg505_out | left_02_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg646_out | left_02_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? right_01_write_out : '0;
  assign left_02_read_write_en = (!(par_done_reg48_out | left_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg78_out | left_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg123_out | left_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg186_out | left_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg270_out | left_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg378_out | left_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg505_out | left_02_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg646_out | left_02_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign top_02_read_in = (!(par_done_reg42_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg68_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg165_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg242_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg342_out | top_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg463_out | top_02_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg600_out | top_02_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? t2_read_data : '0;
  assign top_02_read_write_en = (!(par_done_reg42_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg68_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg165_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg242_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg342_out | top_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg463_out | top_02_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg600_out | top_02_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign pe_02_top = (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? top_02_read_out : '0;
  assign pe_02_left = (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? left_02_read_out : '0;
  assign pe_02_go = (!pe_02_done & (!(par_done_reg62_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg98_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg150_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg221_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg314_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg428_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg559_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg702_out | right_02_write_done & down_02_write_done) & fsm0_out == 32'd21 & !par_reset21_out & go)) ? 1'd1 : '0;
  assign down_01_write_in = (pe_01_done & (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_01_down : '0;
  assign down_01_write_write_en = (pe_01_done & (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign right_01_write_in = (pe_01_done & (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? pe_01_right : '0;
  assign right_01_write_write_en = (pe_01_done & (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign left_01_read_in = (!(par_done_reg29_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg47_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg185_out | left_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg269_out | left_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg377_out | left_01_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg504_out | left_01_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? right_00_write_out : '0;
  assign left_01_read_write_en = (!(par_done_reg29_out | left_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg47_out | left_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg77_out | left_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg122_out | left_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg185_out | left_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg269_out | left_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg377_out | left_01_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg504_out | left_01_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign top_01_read_in = (!(par_done_reg26_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg164_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | top_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg341_out | top_01_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg462_out | top_01_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? t1_read_data : '0;
  assign top_01_read_write_en = (!(par_done_reg26_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg164_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | top_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg341_out | top_01_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg462_out | top_01_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign pe_01_top = (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? top_01_read_out : '0;
  assign pe_01_left = (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? left_01_read_out : '0;
  assign pe_01_go = (!pe_01_done & (!(par_done_reg38_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg61_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg97_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg149_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg220_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg313_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg427_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg558_out | right_01_write_done & down_01_write_done) & fsm0_out == 32'd19 & !par_reset19_out & go)) ? 1'd1 : '0;
  assign down_00_write_in = (pe_00_done & (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_00_down : '0;
  assign down_00_write_write_en = (pe_00_done & (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign right_00_write_in = (pe_00_done & (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? pe_00_right : '0;
  assign right_00_write_write_en = (pe_00_done & (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign left_00_read_in = (!(par_done_reg19_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg28_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg46_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg76_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg121_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg268_out | left_00_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg376_out | left_00_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? l0_read_data : '0;
  assign left_00_read_write_en = (!(par_done_reg19_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg28_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg46_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg76_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg121_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg268_out | left_00_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg376_out | left_00_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign top_00_read_in = (!(par_done_reg18_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg25_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg40_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg66_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | top_00_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg340_out | top_00_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? t0_read_data : '0;
  assign top_00_read_write_en = (!(par_done_reg18_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg25_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg40_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg66_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | top_00_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg340_out | top_00_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign pe_00_top = (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? top_00_read_out : '0;
  assign pe_00_left = (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? left_00_read_out : '0;
  assign pe_00_go = (!pe_00_done & (!(par_done_reg24_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg37_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg60_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg96_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg148_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg219_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg312_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg426_out | right_00_write_done & down_00_write_done) & fsm0_out == 32'd17 & !par_reset17_out & go)) ? 1'd1 : '0;
  assign l7_addr0 = (!(par_done_reg411_out | left_70_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg544_out | left_70_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg689_out | left_70_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg840_out | left_70_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg991_out | left_70_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1136_out | left_70_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1269_out | left_70_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1384_out | left_70_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? l7_idx_out : '0;
  assign l7_add_left = (!(par_done_reg311_out | l7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg425_out | l7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg557_out | l7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg701_out | l7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg851_out | l7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1001_out | l7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1145_out | l7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1277_out | l7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? 4'd1 : '0;
  assign l7_add_right = (!(par_done_reg311_out | l7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg425_out | l7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg557_out | l7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg701_out | l7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg851_out | l7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1001_out | l7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1145_out | l7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1277_out | l7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? l7_idx_out : '0;
  assign l7_idx_in = (!(par_done_reg311_out | l7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg425_out | l7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg557_out | l7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg701_out | l7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg851_out | l7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1001_out | l7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1145_out | l7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1277_out | l7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? l7_add_out : (!(par_done_reg15_out | l7_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l7_idx_write_en = (!(par_done_reg15_out | l7_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg311_out | l7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg425_out | l7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg557_out | l7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg701_out | l7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg851_out | l7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1001_out | l7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1145_out | l7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1277_out | l7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign l6_addr0 = (!(par_done_reg295_out | left_60_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg409_out | left_60_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg541_out | left_60_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg685_out | left_60_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg835_out | left_60_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg985_out | left_60_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1129_out | left_60_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1261_out | left_60_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? l6_idx_out : '0;
  assign l6_add_left = (!(par_done_reg218_out | l6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | l6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg424_out | l6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg556_out | l6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg700_out | l6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg850_out | l6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1000_out | l6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1144_out | l6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? 4'd1 : '0;
  assign l6_add_right = (!(par_done_reg218_out | l6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | l6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg424_out | l6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg556_out | l6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg700_out | l6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg850_out | l6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1000_out | l6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1144_out | l6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? l6_idx_out : '0;
  assign l6_idx_in = (!(par_done_reg218_out | l6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | l6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg424_out | l6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg556_out | l6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg700_out | l6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg850_out | l6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1000_out | l6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1144_out | l6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? l6_add_out : (!(par_done_reg14_out | l6_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l6_idx_write_en = (!(par_done_reg14_out | l6_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg218_out | l6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg310_out | l6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg424_out | l6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg556_out | l6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg700_out | l6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg850_out | l6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg1000_out | l6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1144_out | l6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign l5_addr0 = (!(par_done_reg204_out | left_50_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg293_out | left_50_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg406_out | left_50_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg537_out | left_50_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg680_out | left_50_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg829_out | left_50_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg978_out | left_50_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1121_out | left_50_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? l5_idx_out : '0;
  assign l5_add_left = (!(par_done_reg147_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg309_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg423_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg555_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg699_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg849_out | l5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg999_out | l5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? 4'd1 : '0;
  assign l5_add_right = (!(par_done_reg147_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg309_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg423_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg555_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg699_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg849_out | l5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg999_out | l5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? l5_idx_out : '0;
  assign l5_idx_in = (!(par_done_reg147_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg309_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg423_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg555_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg699_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg849_out | l5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg999_out | l5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? l5_add_out : (!(par_done_reg13_out | l5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l5_idx_write_en = (!(par_done_reg13_out | l5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg147_out | l5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg217_out | l5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg309_out | l5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg423_out | l5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg555_out | l5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg699_out | l5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg849_out | l5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg999_out | l5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign l4_addr0 = (!(par_done_reg135_out | left_40_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg202_out | left_40_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg290_out | left_40_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg402_out | left_40_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg532_out | left_40_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg674_out | left_40_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg822_out | left_40_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg970_out | left_40_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? l4_idx_out : '0;
  assign l4_add_left = (!(par_done_reg95_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg216_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg422_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg554_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg698_out | l4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg848_out | l4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? 4'd1 : '0;
  assign l4_add_right = (!(par_done_reg95_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg216_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg422_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg554_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg698_out | l4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg848_out | l4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? l4_idx_out : '0;
  assign l4_idx_in = (!(par_done_reg95_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg216_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg422_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg554_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg698_out | l4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg848_out | l4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? l4_add_out : (!(par_done_reg12_out | l4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l4_idx_write_en = (!(par_done_reg12_out | l4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg95_out | l4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg146_out | l4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg216_out | l4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg308_out | l4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg422_out | l4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg554_out | l4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg698_out | l4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg848_out | l4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign l3_addr0 = (!(par_done_reg85_out | left_30_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg133_out | left_30_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg199_out | left_30_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg286_out | left_30_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg397_out | left_30_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg526_out | left_30_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg667_out | left_30_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg814_out | left_30_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? l3_idx_out : '0;
  assign l3_add_left = (!(par_done_reg59_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg421_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg553_out | l3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg697_out | l3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 4'd1 : '0;
  assign l3_add_right = (!(par_done_reg59_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg421_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg553_out | l3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg697_out | l3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? l3_idx_out : '0;
  assign l3_idx_in = (!(par_done_reg59_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg421_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg553_out | l3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg697_out | l3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? l3_add_out : (!(par_done_reg11_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l3_idx_write_en = (!(par_done_reg11_out | l3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg59_out | l3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg94_out | l3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg145_out | l3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg215_out | l3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg307_out | l3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg421_out | l3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg553_out | l3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg697_out | l3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign l2_addr0 = (!(par_done_reg51_out | left_20_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg83_out | left_20_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg130_out | left_20_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg195_out | left_20_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg281_out | left_20_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg391_out | left_20_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg519_out | left_20_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg659_out | left_20_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? l2_idx_out : '0;
  assign l2_add_left = (!(par_done_reg36_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg58_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg420_out | l2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg552_out | l2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 4'd1 : '0;
  assign l2_add_right = (!(par_done_reg36_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg58_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg420_out | l2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg552_out | l2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? l2_idx_out : '0;
  assign l2_idx_in = (!(par_done_reg36_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg58_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg420_out | l2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg552_out | l2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? l2_add_out : (!(par_done_reg10_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l2_idx_write_en = (!(par_done_reg10_out | l2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg36_out | l2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg58_out | l2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg93_out | l2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg144_out | l2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg214_out | l2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg306_out | l2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg420_out | l2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg552_out | l2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign l1_addr0 = (!(par_done_reg30_out | left_10_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg49_out | left_10_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg80_out | left_10_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg126_out | left_10_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg190_out | left_10_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg275_out | left_10_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg384_out | left_10_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg511_out | left_10_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? l1_idx_out : '0;
  assign l1_add_left = (!(par_done_reg23_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg35_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg305_out | l1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg419_out | l1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 4'd1 : '0;
  assign l1_add_right = (!(par_done_reg23_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg35_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg305_out | l1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg419_out | l1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? l1_idx_out : '0;
  assign l1_idx_in = (!(par_done_reg23_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg35_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg305_out | l1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg419_out | l1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? l1_add_out : (!(par_done_reg9_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l1_idx_write_en = (!(par_done_reg9_out | l1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg23_out | l1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg35_out | l1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg57_out | l1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg92_out | l1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg143_out | l1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg213_out | l1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg305_out | l1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg419_out | l1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign l0_addr0 = (!(par_done_reg19_out | left_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg28_out | left_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg46_out | left_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg76_out | left_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg121_out | left_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg184_out | left_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg268_out | left_00_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg376_out | left_00_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? l0_idx_out : '0;
  assign l0_add_left = (!(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg21_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg32_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | l0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 4'd1 : '0;
  assign l0_add_right = (!(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg21_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg32_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | l0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? l0_idx_out : '0;
  assign l0_idx_in = (!(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg21_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg32_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | l0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? l0_add_out : (!(par_done_reg8_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign l0_idx_write_en = (!(par_done_reg8_out | l0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg17_out | l0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg21_out | l0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg32_out | l0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg53_out | l0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg87_out | l0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg137_out | l0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg206_out | l0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg297_out | l0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign t7_addr0 = (!(par_done_reg347_out | top_07_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg468_out | top_07_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg605_out | top_07_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg752_out | top_07_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg903_out | top_07_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1052_out | top_07_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1193_out | top_07_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go | !(par_done_reg1320_out | top_07_read_done) & fsm0_out == 32'd30 & !par_reset30_out & go) ? t7_idx_out : '0;
  assign t7_add_left = (!(par_done_reg304_out | t7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg418_out | t7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg551_out | t7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg696_out | t7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg847_out | t7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg998_out | t7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1143_out | t7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1276_out | t7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? 4'd1 : '0;
  assign t7_add_right = (!(par_done_reg304_out | t7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg418_out | t7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg551_out | t7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg696_out | t7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg847_out | t7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg998_out | t7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1143_out | t7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1276_out | t7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? t7_idx_out : '0;
  assign t7_idx_in = (!(par_done_reg304_out | t7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg418_out | t7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg551_out | t7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg696_out | t7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg847_out | t7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg998_out | t7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1143_out | t7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1276_out | t7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? t7_add_out : (!(par_done_reg7_out | t7_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t7_idx_write_en = (!(par_done_reg7_out | t7_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg304_out | t7_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg418_out | t7_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg551_out | t7_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg696_out | t7_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg847_out | t7_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg998_out | t7_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1143_out | t7_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go | !(par_done_reg1276_out | t7_idx_done) & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign t6_addr0 = (!(par_done_reg246_out | top_06_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg346_out | top_06_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg467_out | top_06_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg604_out | top_06_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg751_out | top_06_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg902_out | top_06_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1051_out | top_06_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go | !(par_done_reg1192_out | top_06_read_done) & fsm0_out == 32'd28 & !par_reset28_out & go) ? t6_idx_out : '0;
  assign t6_add_left = (!(par_done_reg212_out | t6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | t6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg417_out | t6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg550_out | t6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg695_out | t6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg846_out | t6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg997_out | t6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1142_out | t6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? 4'd1 : '0;
  assign t6_add_right = (!(par_done_reg212_out | t6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | t6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg417_out | t6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg550_out | t6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg695_out | t6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg846_out | t6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg997_out | t6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1142_out | t6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? t6_idx_out : '0;
  assign t6_idx_in = (!(par_done_reg212_out | t6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | t6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg417_out | t6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg550_out | t6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg695_out | t6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg846_out | t6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg997_out | t6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1142_out | t6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? t6_add_out : (!(par_done_reg6_out | t6_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t6_idx_write_en = (!(par_done_reg6_out | t6_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg212_out | t6_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg303_out | t6_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg417_out | t6_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg550_out | t6_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg695_out | t6_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg846_out | t6_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg997_out | t6_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go | !(par_done_reg1142_out | t6_idx_done) & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign t5_addr0 = (!(par_done_reg168_out | top_05_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg245_out | top_05_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg345_out | top_05_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg466_out | top_05_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg603_out | top_05_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg750_out | top_05_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg901_out | top_05_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go | !(par_done_reg1050_out | top_05_read_done) & fsm0_out == 32'd26 & !par_reset26_out & go) ? t5_idx_out : '0;
  assign t5_add_left = (!(par_done_reg142_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg416_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg549_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg694_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg845_out | t5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg996_out | t5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? 4'd1 : '0;
  assign t5_add_right = (!(par_done_reg142_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg416_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg549_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg694_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg845_out | t5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg996_out | t5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? t5_idx_out : '0;
  assign t5_idx_in = (!(par_done_reg142_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg416_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg549_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg694_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg845_out | t5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg996_out | t5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? t5_add_out : (!(par_done_reg5_out | t5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t5_idx_write_en = (!(par_done_reg5_out | t5_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg142_out | t5_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg211_out | t5_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg302_out | t5_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg416_out | t5_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg549_out | t5_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg694_out | t5_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg845_out | t5_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go | !(par_done_reg996_out | t5_idx_done) & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign t4_addr0 = (!(par_done_reg110_out | top_04_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg167_out | top_04_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg244_out | top_04_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg344_out | top_04_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg465_out | top_04_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg602_out | top_04_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg749_out | top_04_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go | !(par_done_reg900_out | top_04_read_done) & fsm0_out == 32'd24 & !par_reset24_out & go) ? t4_idx_out : '0;
  assign t4_add_left = (!(par_done_reg91_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg415_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg548_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg693_out | t4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg844_out | t4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? 4'd1 : '0;
  assign t4_add_right = (!(par_done_reg91_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg415_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg548_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg693_out | t4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg844_out | t4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? t4_idx_out : '0;
  assign t4_idx_in = (!(par_done_reg91_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg415_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg548_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg693_out | t4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg844_out | t4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? t4_add_out : (!(par_done_reg4_out | t4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t4_idx_write_en = (!(par_done_reg4_out | t4_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg91_out | t4_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg141_out | t4_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg210_out | t4_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg301_out | t4_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg415_out | t4_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg548_out | t4_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg693_out | t4_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go | !(par_done_reg844_out | t4_idx_done) & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign t3_addr0 = (!(par_done_reg69_out | top_03_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg109_out | top_03_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg166_out | top_03_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg243_out | top_03_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg343_out | top_03_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg464_out | top_03_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg601_out | top_03_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go | !(par_done_reg748_out | top_03_read_done) & fsm0_out == 32'd22 & !par_reset22_out & go) ? t3_idx_out : '0;
  assign t3_add_left = (!(par_done_reg56_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg300_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg414_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg547_out | t3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg692_out | t3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 4'd1 : '0;
  assign t3_add_right = (!(par_done_reg56_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg300_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg414_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg547_out | t3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg692_out | t3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? t3_idx_out : '0;
  assign t3_idx_in = (!(par_done_reg56_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg300_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg414_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg547_out | t3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg692_out | t3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? t3_add_out : (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t3_idx_write_en = (!(par_done_reg3_out | t3_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg56_out | t3_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg90_out | t3_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg140_out | t3_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg209_out | t3_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg300_out | t3_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg414_out | t3_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg547_out | t3_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go | !(par_done_reg692_out | t3_idx_done) & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign t2_addr0 = (!(par_done_reg42_out | top_02_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg68_out | top_02_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg108_out | top_02_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg165_out | top_02_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg242_out | top_02_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg342_out | top_02_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg463_out | top_02_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go | !(par_done_reg600_out | top_02_read_done) & fsm0_out == 32'd20 & !par_reset20_out & go) ? t2_idx_out : '0;
  assign t2_add_left = (!(par_done_reg34_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg413_out | t2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg546_out | t2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 4'd1 : '0;
  assign t2_add_right = (!(par_done_reg34_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg413_out | t2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg546_out | t2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? t2_idx_out : '0;
  assign t2_idx_in = (!(par_done_reg34_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg413_out | t2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg546_out | t2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? t2_add_out : (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t2_idx_write_en = (!(par_done_reg2_out | t2_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg34_out | t2_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg55_out | t2_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg89_out | t2_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg139_out | t2_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg208_out | t2_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg299_out | t2_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg413_out | t2_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go | !(par_done_reg546_out | t2_idx_done) & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign t1_addr0 = (!(par_done_reg26_out | top_01_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg41_out | top_01_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg67_out | top_01_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg107_out | top_01_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg164_out | top_01_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg241_out | top_01_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg341_out | top_01_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go | !(par_done_reg462_out | top_01_read_done) & fsm0_out == 32'd18 & !par_reset18_out & go) ? t1_idx_out : '0;
  assign t1_add_left = (!(par_done_reg22_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | t1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg412_out | t1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 4'd1 : '0;
  assign t1_add_right = (!(par_done_reg22_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | t1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg412_out | t1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? t1_idx_out : '0;
  assign t1_idx_in = (!(par_done_reg22_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | t1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg412_out | t1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? t1_add_out : (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t1_idx_write_en = (!(par_done_reg1_out | t1_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg22_out | t1_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg33_out | t1_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg54_out | t1_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg88_out | t1_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg138_out | t1_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg207_out | t1_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg298_out | t1_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go | !(par_done_reg412_out | t1_idx_done) & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign t0_addr0 = (!(par_done_reg18_out | top_00_read_done) & fsm0_out == 32'd2 & !par_reset2_out & go | !(par_done_reg25_out | top_00_read_done) & fsm0_out == 32'd4 & !par_reset4_out & go | !(par_done_reg40_out | top_00_read_done) & fsm0_out == 32'd6 & !par_reset6_out & go | !(par_done_reg66_out | top_00_read_done) & fsm0_out == 32'd8 & !par_reset8_out & go | !(par_done_reg106_out | top_00_read_done) & fsm0_out == 32'd10 & !par_reset10_out & go | !(par_done_reg163_out | top_00_read_done) & fsm0_out == 32'd12 & !par_reset12_out & go | !(par_done_reg240_out | top_00_read_done) & fsm0_out == 32'd14 & !par_reset14_out & go | !(par_done_reg340_out | top_00_read_done) & fsm0_out == 32'd16 & !par_reset16_out & go) ? t0_idx_out : '0;
  assign t0_add_left = (!(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg20_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | t0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 4'd1 : '0;
  assign t0_add_right = (!(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg20_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | t0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? t0_idx_out : '0;
  assign t0_idx_in = (!(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg20_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | t0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? t0_add_out : (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go) ? 4'd15 : '0;
  assign t0_idx_write_en = (!(par_done_reg0_out | t0_idx_done) & fsm0_out == 32'd0 & !par_reset0_out & go | !(par_done_reg16_out | t0_idx_done) & fsm0_out == 32'd1 & !par_reset1_out & go | !(par_done_reg20_out | t0_idx_done) & fsm0_out == 32'd3 & !par_reset3_out & go | !(par_done_reg31_out | t0_idx_done) & fsm0_out == 32'd5 & !par_reset5_out & go | !(par_done_reg52_out | t0_idx_done) & fsm0_out == 32'd7 & !par_reset7_out & go | !(par_done_reg86_out | t0_idx_done) & fsm0_out == 32'd9 & !par_reset9_out & go | !(par_done_reg136_out | t0_idx_done) & fsm0_out == 32'd11 & !par_reset11_out & go | !(par_done_reg205_out | t0_idx_done) & fsm0_out == 32'd13 & !par_reset13_out & go | !(par_done_reg296_out | t0_idx_done) & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_reset0_in = par_reset0_out ? 1'd0 : (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & par_done_reg8_out & par_done_reg9_out & par_done_reg10_out & par_done_reg11_out & par_done_reg12_out & par_done_reg13_out & par_done_reg14_out & par_done_reg15_out & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_reset0_write_en = (par_done_reg0_out & par_done_reg1_out & par_done_reg2_out & par_done_reg3_out & par_done_reg4_out & par_done_reg5_out & par_done_reg6_out & par_done_reg7_out & par_done_reg8_out & par_done_reg9_out & par_done_reg10_out & par_done_reg11_out & par_done_reg12_out & par_done_reg13_out & par_done_reg14_out & par_done_reg15_out & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg0_in = par_reset0_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg0_write_en = (t0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg1_in = par_reset0_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg1_write_en = (t1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg2_in = par_reset0_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg2_write_en = (t2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg3_in = par_reset0_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg3_write_en = (t3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg4_in = par_reset0_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg4_write_en = (t4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg5_in = par_reset0_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg5_write_en = (t5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg6_in = par_reset0_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg6_write_en = (t6_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg7_in = par_reset0_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg7_write_en = (t7_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg8_in = par_reset0_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg8_write_en = (l0_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg9_in = par_reset0_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg9_write_en = (l1_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg10_in = par_reset0_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg10_write_en = (l2_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg11_in = par_reset0_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg11_write_en = (l3_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg12_in = par_reset0_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg12_write_en = (l4_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg13_in = par_reset0_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg13_write_en = (l5_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg14_in = par_reset0_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg14_write_en = (l6_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_done_reg15_in = par_reset0_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go) ? 1'd1 : '0;
  assign par_done_reg15_write_en = (l7_idx_done & fsm0_out == 32'd0 & !par_reset0_out & go | par_reset0_out) ? 1'd1 : '0;
  assign par_reset1_in = par_reset1_out ? 1'd0 : (par_done_reg16_out & par_done_reg17_out & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_reset1_write_en = (par_done_reg16_out & par_done_reg17_out & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg16_in = par_reset1_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg16_write_en = (t0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_done_reg17_in = par_reset1_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go) ? 1'd1 : '0;
  assign par_done_reg17_write_en = (l0_idx_done & fsm0_out == 32'd1 & !par_reset1_out & go | par_reset1_out) ? 1'd1 : '0;
  assign par_reset2_in = par_reset2_out ? 1'd0 : (par_done_reg18_out & par_done_reg19_out & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_reset2_write_en = (par_done_reg18_out & par_done_reg19_out & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg18_in = par_reset2_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg18_write_en = (top_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_done_reg19_in = par_reset2_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go) ? 1'd1 : '0;
  assign par_done_reg19_write_en = (left_00_read_done & fsm0_out == 32'd2 & !par_reset2_out & go | par_reset2_out) ? 1'd1 : '0;
  assign par_reset3_in = par_reset3_out ? 1'd0 : (par_done_reg20_out & par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_reset3_write_en = (par_done_reg20_out & par_done_reg21_out & par_done_reg22_out & par_done_reg23_out & par_done_reg24_out & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg20_in = par_reset3_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg20_write_en = (t0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg21_in = par_reset3_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg21_write_en = (l0_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg22_in = par_reset3_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg22_write_en = (t1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg23_in = par_reset3_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg23_write_en = (l1_idx_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_done_reg24_in = par_reset3_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go) ? 1'd1 : '0;
  assign par_done_reg24_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd3 & !par_reset3_out & go | par_reset3_out) ? 1'd1 : '0;
  assign par_reset4_in = par_reset4_out ? 1'd0 : (par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_reset4_write_en = (par_done_reg25_out & par_done_reg26_out & par_done_reg27_out & par_done_reg28_out & par_done_reg29_out & par_done_reg30_out & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg25_in = par_reset4_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg25_write_en = (top_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg26_in = par_reset4_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg26_write_en = (top_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg27_in = par_reset4_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg27_write_en = (top_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg28_in = par_reset4_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg28_write_en = (left_00_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg29_in = par_reset4_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg29_write_en = (left_01_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_done_reg30_in = par_reset4_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go) ? 1'd1 : '0;
  assign par_done_reg30_write_en = (left_10_read_done & fsm0_out == 32'd4 & !par_reset4_out & go | par_reset4_out) ? 1'd1 : '0;
  assign par_reset5_in = par_reset5_out ? 1'd0 : (par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_reset5_write_en = (par_done_reg31_out & par_done_reg32_out & par_done_reg33_out & par_done_reg34_out & par_done_reg35_out & par_done_reg36_out & par_done_reg37_out & par_done_reg38_out & par_done_reg39_out & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg31_in = par_reset5_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg31_write_en = (t0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg32_in = par_reset5_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg32_write_en = (l0_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg33_in = par_reset5_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg33_write_en = (t1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg34_in = par_reset5_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg34_write_en = (t2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg35_in = par_reset5_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg35_write_en = (l1_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg36_in = par_reset5_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg36_write_en = (l2_idx_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg37_in = par_reset5_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg37_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg38_in = par_reset5_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg38_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_done_reg39_in = par_reset5_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go) ? 1'd1 : '0;
  assign par_done_reg39_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd5 & !par_reset5_out & go | par_reset5_out) ? 1'd1 : '0;
  assign par_reset6_in = par_reset6_out ? 1'd0 : (par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_reset6_write_en = (par_done_reg40_out & par_done_reg41_out & par_done_reg42_out & par_done_reg43_out & par_done_reg44_out & par_done_reg45_out & par_done_reg46_out & par_done_reg47_out & par_done_reg48_out & par_done_reg49_out & par_done_reg50_out & par_done_reg51_out & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg40_in = par_reset6_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg40_write_en = (top_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg41_in = par_reset6_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg41_write_en = (top_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg42_in = par_reset6_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg42_write_en = (top_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg43_in = par_reset6_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg43_write_en = (top_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg44_in = par_reset6_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg44_write_en = (top_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg45_in = par_reset6_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg45_write_en = (top_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg46_in = par_reset6_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg46_write_en = (left_00_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg47_in = par_reset6_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg47_write_en = (left_01_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg48_in = par_reset6_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg48_write_en = (left_02_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg49_in = par_reset6_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg49_write_en = (left_10_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg50_in = par_reset6_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg50_write_en = (left_11_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_done_reg51_in = par_reset6_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go) ? 1'd1 : '0;
  assign par_done_reg51_write_en = (left_20_read_done & fsm0_out == 32'd6 & !par_reset6_out & go | par_reset6_out) ? 1'd1 : '0;
  assign par_reset7_in = par_reset7_out ? 1'd0 : (par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_reset7_write_en = (par_done_reg52_out & par_done_reg53_out & par_done_reg54_out & par_done_reg55_out & par_done_reg56_out & par_done_reg57_out & par_done_reg58_out & par_done_reg59_out & par_done_reg60_out & par_done_reg61_out & par_done_reg62_out & par_done_reg63_out & par_done_reg64_out & par_done_reg65_out & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg52_in = par_reset7_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg52_write_en = (t0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg53_in = par_reset7_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg53_write_en = (l0_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg54_in = par_reset7_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg54_write_en = (t1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg55_in = par_reset7_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg55_write_en = (t2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg56_in = par_reset7_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg56_write_en = (t3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg57_in = par_reset7_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg57_write_en = (l1_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg58_in = par_reset7_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg58_write_en = (l2_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg59_in = par_reset7_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg59_write_en = (l3_idx_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg60_in = par_reset7_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg60_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg61_in = par_reset7_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg61_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg62_in = par_reset7_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg62_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg63_in = par_reset7_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg63_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg64_in = par_reset7_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg64_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_done_reg65_in = par_reset7_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go) ? 1'd1 : '0;
  assign par_done_reg65_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd7 & !par_reset7_out & go | par_reset7_out) ? 1'd1 : '0;
  assign par_reset8_in = par_reset8_out ? 1'd0 : (par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_reset8_write_en = (par_done_reg66_out & par_done_reg67_out & par_done_reg68_out & par_done_reg69_out & par_done_reg70_out & par_done_reg71_out & par_done_reg72_out & par_done_reg73_out & par_done_reg74_out & par_done_reg75_out & par_done_reg76_out & par_done_reg77_out & par_done_reg78_out & par_done_reg79_out & par_done_reg80_out & par_done_reg81_out & par_done_reg82_out & par_done_reg83_out & par_done_reg84_out & par_done_reg85_out & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg66_in = par_reset8_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg66_write_en = (top_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg67_in = par_reset8_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg67_write_en = (top_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg68_in = par_reset8_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg68_write_en = (top_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg69_in = par_reset8_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg69_write_en = (top_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg70_in = par_reset8_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg70_write_en = (top_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg71_in = par_reset8_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg71_write_en = (top_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg72_in = par_reset8_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg72_write_en = (top_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg73_in = par_reset8_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg73_write_en = (top_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg74_in = par_reset8_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg74_write_en = (top_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg75_in = par_reset8_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg75_write_en = (top_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg76_in = par_reset8_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg76_write_en = (left_00_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg77_in = par_reset8_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg77_write_en = (left_01_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg78_in = par_reset8_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg78_write_en = (left_02_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg79_in = par_reset8_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg79_write_en = (left_03_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg80_in = par_reset8_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg80_write_en = (left_10_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg81_in = par_reset8_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg81_write_en = (left_11_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg82_in = par_reset8_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg82_write_en = (left_12_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg83_in = par_reset8_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg83_write_en = (left_20_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg84_in = par_reset8_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg84_write_en = (left_21_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_done_reg85_in = par_reset8_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go) ? 1'd1 : '0;
  assign par_done_reg85_write_en = (left_30_read_done & fsm0_out == 32'd8 & !par_reset8_out & go | par_reset8_out) ? 1'd1 : '0;
  assign par_reset9_in = par_reset9_out ? 1'd0 : (par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_reset9_write_en = (par_done_reg86_out & par_done_reg87_out & par_done_reg88_out & par_done_reg89_out & par_done_reg90_out & par_done_reg91_out & par_done_reg92_out & par_done_reg93_out & par_done_reg94_out & par_done_reg95_out & par_done_reg96_out & par_done_reg97_out & par_done_reg98_out & par_done_reg99_out & par_done_reg100_out & par_done_reg101_out & par_done_reg102_out & par_done_reg103_out & par_done_reg104_out & par_done_reg105_out & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg86_in = par_reset9_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg86_write_en = (t0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg87_in = par_reset9_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg87_write_en = (l0_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg88_in = par_reset9_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg88_write_en = (t1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg89_in = par_reset9_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg89_write_en = (t2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg90_in = par_reset9_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg90_write_en = (t3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg91_in = par_reset9_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg91_write_en = (t4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg92_in = par_reset9_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg92_write_en = (l1_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg93_in = par_reset9_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg93_write_en = (l2_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg94_in = par_reset9_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg94_write_en = (l3_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg95_in = par_reset9_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg95_write_en = (l4_idx_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg96_in = par_reset9_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg96_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg97_in = par_reset9_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg97_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg98_in = par_reset9_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg98_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg99_in = par_reset9_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg99_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg100_in = par_reset9_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg100_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg101_in = par_reset9_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg101_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg102_in = par_reset9_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg102_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg103_in = par_reset9_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg103_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg104_in = par_reset9_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg104_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_done_reg105_in = par_reset9_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go) ? 1'd1 : '0;
  assign par_done_reg105_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd9 & !par_reset9_out & go | par_reset9_out) ? 1'd1 : '0;
  assign par_reset10_in = par_reset10_out ? 1'd0 : (par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & par_done_reg130_out & par_done_reg131_out & par_done_reg132_out & par_done_reg133_out & par_done_reg134_out & par_done_reg135_out & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_reset10_write_en = (par_done_reg106_out & par_done_reg107_out & par_done_reg108_out & par_done_reg109_out & par_done_reg110_out & par_done_reg111_out & par_done_reg112_out & par_done_reg113_out & par_done_reg114_out & par_done_reg115_out & par_done_reg116_out & par_done_reg117_out & par_done_reg118_out & par_done_reg119_out & par_done_reg120_out & par_done_reg121_out & par_done_reg122_out & par_done_reg123_out & par_done_reg124_out & par_done_reg125_out & par_done_reg126_out & par_done_reg127_out & par_done_reg128_out & par_done_reg129_out & par_done_reg130_out & par_done_reg131_out & par_done_reg132_out & par_done_reg133_out & par_done_reg134_out & par_done_reg135_out & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg106_in = par_reset10_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg106_write_en = (top_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg107_in = par_reset10_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg107_write_en = (top_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg108_in = par_reset10_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg108_write_en = (top_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg109_in = par_reset10_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg109_write_en = (top_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg110_in = par_reset10_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg110_write_en = (top_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg111_in = par_reset10_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg111_write_en = (top_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg112_in = par_reset10_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg112_write_en = (top_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg113_in = par_reset10_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg113_write_en = (top_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg114_in = par_reset10_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg114_write_en = (top_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg115_in = par_reset10_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg115_write_en = (top_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg116_in = par_reset10_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg116_write_en = (top_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg117_in = par_reset10_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg117_write_en = (top_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg118_in = par_reset10_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg118_write_en = (top_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg119_in = par_reset10_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg119_write_en = (top_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg120_in = par_reset10_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg120_write_en = (top_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg121_in = par_reset10_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg121_write_en = (left_00_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg122_in = par_reset10_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg122_write_en = (left_01_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg123_in = par_reset10_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg123_write_en = (left_02_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg124_in = par_reset10_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg124_write_en = (left_03_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg125_in = par_reset10_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg125_write_en = (left_04_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg126_in = par_reset10_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg126_write_en = (left_10_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg127_in = par_reset10_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg127_write_en = (left_11_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg128_in = par_reset10_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg128_write_en = (left_12_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg129_in = par_reset10_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg129_write_en = (left_13_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg130_in = par_reset10_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg130_write_en = (left_20_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg131_in = par_reset10_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg131_write_en = (left_21_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg132_in = par_reset10_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg132_write_en = (left_22_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg133_in = par_reset10_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg133_write_en = (left_30_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg134_in = par_reset10_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg134_write_en = (left_31_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_done_reg135_in = par_reset10_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go) ? 1'd1 : '0;
  assign par_done_reg135_write_en = (left_40_read_done & fsm0_out == 32'd10 & !par_reset10_out & go | par_reset10_out) ? 1'd1 : '0;
  assign par_reset11_in = par_reset11_out ? 1'd0 : (par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & par_done_reg158_out & par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_reset11_write_en = (par_done_reg136_out & par_done_reg137_out & par_done_reg138_out & par_done_reg139_out & par_done_reg140_out & par_done_reg141_out & par_done_reg142_out & par_done_reg143_out & par_done_reg144_out & par_done_reg145_out & par_done_reg146_out & par_done_reg147_out & par_done_reg148_out & par_done_reg149_out & par_done_reg150_out & par_done_reg151_out & par_done_reg152_out & par_done_reg153_out & par_done_reg154_out & par_done_reg155_out & par_done_reg156_out & par_done_reg157_out & par_done_reg158_out & par_done_reg159_out & par_done_reg160_out & par_done_reg161_out & par_done_reg162_out & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg136_in = par_reset11_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg136_write_en = (t0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg137_in = par_reset11_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg137_write_en = (l0_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg138_in = par_reset11_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg138_write_en = (t1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg139_in = par_reset11_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg139_write_en = (t2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg140_in = par_reset11_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg140_write_en = (t3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg141_in = par_reset11_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg141_write_en = (t4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg142_in = par_reset11_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg142_write_en = (t5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg143_in = par_reset11_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg143_write_en = (l1_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg144_in = par_reset11_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg144_write_en = (l2_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg145_in = par_reset11_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg145_write_en = (l3_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg146_in = par_reset11_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg146_write_en = (l4_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg147_in = par_reset11_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg147_write_en = (l5_idx_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg148_in = par_reset11_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg148_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg149_in = par_reset11_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg149_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg150_in = par_reset11_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg150_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg151_in = par_reset11_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg151_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg152_in = par_reset11_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg152_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg153_in = par_reset11_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg153_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg154_in = par_reset11_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg154_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg155_in = par_reset11_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg155_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg156_in = par_reset11_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg156_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg157_in = par_reset11_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg157_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg158_in = par_reset11_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg158_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg159_in = par_reset11_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg159_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg160_in = par_reset11_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg160_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg161_in = par_reset11_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg161_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_done_reg162_in = par_reset11_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd11 & !par_reset11_out & go) ? 1'd1 : '0;
  assign par_done_reg162_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd11 & !par_reset11_out & go | par_reset11_out) ? 1'd1 : '0;
  assign par_reset12_in = par_reset12_out ? 1'd0 : (par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & par_done_reg201_out & par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_reset12_write_en = (par_done_reg163_out & par_done_reg164_out & par_done_reg165_out & par_done_reg166_out & par_done_reg167_out & par_done_reg168_out & par_done_reg169_out & par_done_reg170_out & par_done_reg171_out & par_done_reg172_out & par_done_reg173_out & par_done_reg174_out & par_done_reg175_out & par_done_reg176_out & par_done_reg177_out & par_done_reg178_out & par_done_reg179_out & par_done_reg180_out & par_done_reg181_out & par_done_reg182_out & par_done_reg183_out & par_done_reg184_out & par_done_reg185_out & par_done_reg186_out & par_done_reg187_out & par_done_reg188_out & par_done_reg189_out & par_done_reg190_out & par_done_reg191_out & par_done_reg192_out & par_done_reg193_out & par_done_reg194_out & par_done_reg195_out & par_done_reg196_out & par_done_reg197_out & par_done_reg198_out & par_done_reg199_out & par_done_reg200_out & par_done_reg201_out & par_done_reg202_out & par_done_reg203_out & par_done_reg204_out & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg163_in = par_reset12_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg163_write_en = (top_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg164_in = par_reset12_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg164_write_en = (top_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg165_in = par_reset12_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg165_write_en = (top_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg166_in = par_reset12_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg166_write_en = (top_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg167_in = par_reset12_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg167_write_en = (top_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg168_in = par_reset12_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg168_write_en = (top_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg169_in = par_reset12_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg169_write_en = (top_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg170_in = par_reset12_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg170_write_en = (top_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg171_in = par_reset12_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg171_write_en = (top_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg172_in = par_reset12_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg172_write_en = (top_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg173_in = par_reset12_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg173_write_en = (top_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg174_in = par_reset12_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg174_write_en = (top_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg175_in = par_reset12_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg175_write_en = (top_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg176_in = par_reset12_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg176_write_en = (top_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg177_in = par_reset12_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg177_write_en = (top_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg178_in = par_reset12_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg178_write_en = (top_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg179_in = par_reset12_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg179_write_en = (top_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg180_in = par_reset12_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg180_write_en = (top_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg181_in = par_reset12_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg181_write_en = (top_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg182_in = par_reset12_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg182_write_en = (top_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg183_in = par_reset12_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg183_write_en = (top_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg184_in = par_reset12_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg184_write_en = (left_00_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg185_in = par_reset12_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg185_write_en = (left_01_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg186_in = par_reset12_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg186_write_en = (left_02_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg187_in = par_reset12_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg187_write_en = (left_03_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg188_in = par_reset12_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg188_write_en = (left_04_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg189_in = par_reset12_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg189_write_en = (left_05_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg190_in = par_reset12_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg190_write_en = (left_10_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg191_in = par_reset12_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg191_write_en = (left_11_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg192_in = par_reset12_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg192_write_en = (left_12_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg193_in = par_reset12_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg193_write_en = (left_13_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg194_in = par_reset12_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg194_write_en = (left_14_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg195_in = par_reset12_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg195_write_en = (left_20_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg196_in = par_reset12_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg196_write_en = (left_21_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg197_in = par_reset12_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg197_write_en = (left_22_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg198_in = par_reset12_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg198_write_en = (left_23_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg199_in = par_reset12_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg199_write_en = (left_30_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg200_in = par_reset12_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg200_write_en = (left_31_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg201_in = par_reset12_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg201_write_en = (left_32_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg202_in = par_reset12_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg202_write_en = (left_40_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg203_in = par_reset12_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg203_write_en = (left_41_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_done_reg204_in = par_reset12_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go) ? 1'd1 : '0;
  assign par_done_reg204_write_en = (left_50_read_done & fsm0_out == 32'd12 & !par_reset12_out & go | par_reset12_out) ? 1'd1 : '0;
  assign par_reset13_in = par_reset13_out ? 1'd0 : (par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & par_done_reg213_out & par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & par_done_reg229_out & par_done_reg230_out & par_done_reg231_out & par_done_reg232_out & par_done_reg233_out & par_done_reg234_out & par_done_reg235_out & par_done_reg236_out & par_done_reg237_out & par_done_reg238_out & par_done_reg239_out & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_reset13_write_en = (par_done_reg205_out & par_done_reg206_out & par_done_reg207_out & par_done_reg208_out & par_done_reg209_out & par_done_reg210_out & par_done_reg211_out & par_done_reg212_out & par_done_reg213_out & par_done_reg214_out & par_done_reg215_out & par_done_reg216_out & par_done_reg217_out & par_done_reg218_out & par_done_reg219_out & par_done_reg220_out & par_done_reg221_out & par_done_reg222_out & par_done_reg223_out & par_done_reg224_out & par_done_reg225_out & par_done_reg226_out & par_done_reg227_out & par_done_reg228_out & par_done_reg229_out & par_done_reg230_out & par_done_reg231_out & par_done_reg232_out & par_done_reg233_out & par_done_reg234_out & par_done_reg235_out & par_done_reg236_out & par_done_reg237_out & par_done_reg238_out & par_done_reg239_out & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg205_in = par_reset13_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg205_write_en = (t0_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg206_in = par_reset13_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg206_write_en = (l0_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg207_in = par_reset13_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg207_write_en = (t1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg208_in = par_reset13_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg208_write_en = (t2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg209_in = par_reset13_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg209_write_en = (t3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg210_in = par_reset13_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg210_write_en = (t4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg211_in = par_reset13_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg211_write_en = (t5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg212_in = par_reset13_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg212_write_en = (t6_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg213_in = par_reset13_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg213_write_en = (l1_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg214_in = par_reset13_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg214_write_en = (l2_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg215_in = par_reset13_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg215_write_en = (l3_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg216_in = par_reset13_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg216_write_en = (l4_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg217_in = par_reset13_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg217_write_en = (l5_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg218_in = par_reset13_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg218_write_en = (l6_idx_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg219_in = par_reset13_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg219_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg220_in = par_reset13_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg220_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg221_in = par_reset13_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg221_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg222_in = par_reset13_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg222_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg223_in = par_reset13_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg223_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg224_in = par_reset13_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg224_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg225_in = par_reset13_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg225_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg226_in = par_reset13_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg226_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg227_in = par_reset13_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg227_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg228_in = par_reset13_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg228_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg229_in = par_reset13_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg229_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg230_in = par_reset13_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg230_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg231_in = par_reset13_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg231_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg232_in = par_reset13_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg232_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg233_in = par_reset13_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg233_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg234_in = par_reset13_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg234_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg235_in = par_reset13_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg235_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg236_in = par_reset13_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg236_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg237_in = par_reset13_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg237_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg238_in = par_reset13_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg238_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_done_reg239_in = par_reset13_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd13 & !par_reset13_out & go) ? 1'd1 : '0;
  assign par_done_reg239_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd13 & !par_reset13_out & go | par_reset13_out) ? 1'd1 : '0;
  assign par_reset14_in = par_reset14_out ? 1'd0 : (par_done_reg240_out & par_done_reg241_out & par_done_reg242_out & par_done_reg243_out & par_done_reg244_out & par_done_reg245_out & par_done_reg246_out & par_done_reg247_out & par_done_reg248_out & par_done_reg249_out & par_done_reg250_out & par_done_reg251_out & par_done_reg252_out & par_done_reg253_out & par_done_reg254_out & par_done_reg255_out & par_done_reg256_out & par_done_reg257_out & par_done_reg258_out & par_done_reg259_out & par_done_reg260_out & par_done_reg261_out & par_done_reg262_out & par_done_reg263_out & par_done_reg264_out & par_done_reg265_out & par_done_reg266_out & par_done_reg267_out & par_done_reg268_out & par_done_reg269_out & par_done_reg270_out & par_done_reg271_out & par_done_reg272_out & par_done_reg273_out & par_done_reg274_out & par_done_reg275_out & par_done_reg276_out & par_done_reg277_out & par_done_reg278_out & par_done_reg279_out & par_done_reg280_out & par_done_reg281_out & par_done_reg282_out & par_done_reg283_out & par_done_reg284_out & par_done_reg285_out & par_done_reg286_out & par_done_reg287_out & par_done_reg288_out & par_done_reg289_out & par_done_reg290_out & par_done_reg291_out & par_done_reg292_out & par_done_reg293_out & par_done_reg294_out & par_done_reg295_out & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_reset14_write_en = (par_done_reg240_out & par_done_reg241_out & par_done_reg242_out & par_done_reg243_out & par_done_reg244_out & par_done_reg245_out & par_done_reg246_out & par_done_reg247_out & par_done_reg248_out & par_done_reg249_out & par_done_reg250_out & par_done_reg251_out & par_done_reg252_out & par_done_reg253_out & par_done_reg254_out & par_done_reg255_out & par_done_reg256_out & par_done_reg257_out & par_done_reg258_out & par_done_reg259_out & par_done_reg260_out & par_done_reg261_out & par_done_reg262_out & par_done_reg263_out & par_done_reg264_out & par_done_reg265_out & par_done_reg266_out & par_done_reg267_out & par_done_reg268_out & par_done_reg269_out & par_done_reg270_out & par_done_reg271_out & par_done_reg272_out & par_done_reg273_out & par_done_reg274_out & par_done_reg275_out & par_done_reg276_out & par_done_reg277_out & par_done_reg278_out & par_done_reg279_out & par_done_reg280_out & par_done_reg281_out & par_done_reg282_out & par_done_reg283_out & par_done_reg284_out & par_done_reg285_out & par_done_reg286_out & par_done_reg287_out & par_done_reg288_out & par_done_reg289_out & par_done_reg290_out & par_done_reg291_out & par_done_reg292_out & par_done_reg293_out & par_done_reg294_out & par_done_reg295_out & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg240_in = par_reset14_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg240_write_en = (top_00_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg241_in = par_reset14_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg241_write_en = (top_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg242_in = par_reset14_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg242_write_en = (top_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg243_in = par_reset14_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg243_write_en = (top_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg244_in = par_reset14_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg244_write_en = (top_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg245_in = par_reset14_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg245_write_en = (top_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg246_in = par_reset14_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg246_write_en = (top_06_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg247_in = par_reset14_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg247_write_en = (top_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg248_in = par_reset14_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg248_write_en = (top_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg249_in = par_reset14_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg249_write_en = (top_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg250_in = par_reset14_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg250_write_en = (top_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg251_in = par_reset14_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg251_write_en = (top_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg252_in = par_reset14_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg252_write_en = (top_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg253_in = par_reset14_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg253_write_en = (top_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg254_in = par_reset14_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg254_write_en = (top_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg255_in = par_reset14_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg255_write_en = (top_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg256_in = par_reset14_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg256_write_en = (top_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg257_in = par_reset14_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg257_write_en = (top_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg258_in = par_reset14_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg258_write_en = (top_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg259_in = par_reset14_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg259_write_en = (top_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg260_in = par_reset14_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg260_write_en = (top_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg261_in = par_reset14_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg261_write_en = (top_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg262_in = par_reset14_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg262_write_en = (top_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg263_in = par_reset14_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg263_write_en = (top_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg264_in = par_reset14_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg264_write_en = (top_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg265_in = par_reset14_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg265_write_en = (top_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg266_in = par_reset14_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg266_write_en = (top_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg267_in = par_reset14_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg267_write_en = (top_60_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg268_in = par_reset14_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg268_write_en = (left_00_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg269_in = par_reset14_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg269_write_en = (left_01_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg270_in = par_reset14_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg270_write_en = (left_02_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg271_in = par_reset14_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg271_write_en = (left_03_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg272_in = par_reset14_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg272_write_en = (left_04_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg273_in = par_reset14_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg273_write_en = (left_05_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg274_in = par_reset14_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg274_write_en = (left_06_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg275_in = par_reset14_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg275_write_en = (left_10_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg276_in = par_reset14_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg276_write_en = (left_11_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg277_in = par_reset14_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg277_write_en = (left_12_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg278_in = par_reset14_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg278_write_en = (left_13_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg279_in = par_reset14_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg279_write_en = (left_14_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg280_in = par_reset14_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg280_write_en = (left_15_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg281_in = par_reset14_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg281_write_en = (left_20_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg282_in = par_reset14_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg282_write_en = (left_21_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg283_in = par_reset14_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg283_write_en = (left_22_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg284_in = par_reset14_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg284_write_en = (left_23_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg285_in = par_reset14_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg285_write_en = (left_24_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg286_in = par_reset14_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg286_write_en = (left_30_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg287_in = par_reset14_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg287_write_en = (left_31_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg288_in = par_reset14_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg288_write_en = (left_32_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg289_in = par_reset14_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg289_write_en = (left_33_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg290_in = par_reset14_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg290_write_en = (left_40_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg291_in = par_reset14_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg291_write_en = (left_41_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg292_in = par_reset14_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg292_write_en = (left_42_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg293_in = par_reset14_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg293_write_en = (left_50_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg294_in = par_reset14_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg294_write_en = (left_51_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_done_reg295_in = par_reset14_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd14 & !par_reset14_out & go) ? 1'd1 : '0;
  assign par_done_reg295_write_en = (left_60_read_done & fsm0_out == 32'd14 & !par_reset14_out & go | par_reset14_out) ? 1'd1 : '0;
  assign par_reset15_in = par_reset15_out ? 1'd0 : (par_done_reg296_out & par_done_reg297_out & par_done_reg298_out & par_done_reg299_out & par_done_reg300_out & par_done_reg301_out & par_done_reg302_out & par_done_reg303_out & par_done_reg304_out & par_done_reg305_out & par_done_reg306_out & par_done_reg307_out & par_done_reg308_out & par_done_reg309_out & par_done_reg310_out & par_done_reg311_out & par_done_reg312_out & par_done_reg313_out & par_done_reg314_out & par_done_reg315_out & par_done_reg316_out & par_done_reg317_out & par_done_reg318_out & par_done_reg319_out & par_done_reg320_out & par_done_reg321_out & par_done_reg322_out & par_done_reg323_out & par_done_reg324_out & par_done_reg325_out & par_done_reg326_out & par_done_reg327_out & par_done_reg328_out & par_done_reg329_out & par_done_reg330_out & par_done_reg331_out & par_done_reg332_out & par_done_reg333_out & par_done_reg334_out & par_done_reg335_out & par_done_reg336_out & par_done_reg337_out & par_done_reg338_out & par_done_reg339_out & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_reset15_write_en = (par_done_reg296_out & par_done_reg297_out & par_done_reg298_out & par_done_reg299_out & par_done_reg300_out & par_done_reg301_out & par_done_reg302_out & par_done_reg303_out & par_done_reg304_out & par_done_reg305_out & par_done_reg306_out & par_done_reg307_out & par_done_reg308_out & par_done_reg309_out & par_done_reg310_out & par_done_reg311_out & par_done_reg312_out & par_done_reg313_out & par_done_reg314_out & par_done_reg315_out & par_done_reg316_out & par_done_reg317_out & par_done_reg318_out & par_done_reg319_out & par_done_reg320_out & par_done_reg321_out & par_done_reg322_out & par_done_reg323_out & par_done_reg324_out & par_done_reg325_out & par_done_reg326_out & par_done_reg327_out & par_done_reg328_out & par_done_reg329_out & par_done_reg330_out & par_done_reg331_out & par_done_reg332_out & par_done_reg333_out & par_done_reg334_out & par_done_reg335_out & par_done_reg336_out & par_done_reg337_out & par_done_reg338_out & par_done_reg339_out & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg296_in = par_reset15_out ? 1'd0 : (t0_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg296_write_en = (t0_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg297_in = par_reset15_out ? 1'd0 : (l0_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg297_write_en = (l0_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg298_in = par_reset15_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg298_write_en = (t1_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg299_in = par_reset15_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg299_write_en = (t2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg300_in = par_reset15_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg300_write_en = (t3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg301_in = par_reset15_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg301_write_en = (t4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg302_in = par_reset15_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg302_write_en = (t5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg303_in = par_reset15_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg303_write_en = (t6_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg304_in = par_reset15_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg304_write_en = (t7_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg305_in = par_reset15_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg305_write_en = (l1_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg306_in = par_reset15_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg306_write_en = (l2_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg307_in = par_reset15_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg307_write_en = (l3_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg308_in = par_reset15_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg308_write_en = (l4_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg309_in = par_reset15_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg309_write_en = (l5_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg310_in = par_reset15_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg310_write_en = (l6_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg311_in = par_reset15_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg311_write_en = (l7_idx_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg312_in = par_reset15_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg312_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg313_in = par_reset15_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg313_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg314_in = par_reset15_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg314_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg315_in = par_reset15_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg315_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg316_in = par_reset15_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg316_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg317_in = par_reset15_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg317_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg318_in = par_reset15_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg318_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg319_in = par_reset15_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg319_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg320_in = par_reset15_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg320_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg321_in = par_reset15_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg321_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg322_in = par_reset15_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg322_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg323_in = par_reset15_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg323_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg324_in = par_reset15_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg324_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg325_in = par_reset15_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg325_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg326_in = par_reset15_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg326_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg327_in = par_reset15_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg327_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg328_in = par_reset15_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg328_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg329_in = par_reset15_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg329_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg330_in = par_reset15_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg330_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg331_in = par_reset15_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg331_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg332_in = par_reset15_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg332_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg333_in = par_reset15_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg333_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg334_in = par_reset15_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg334_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg335_in = par_reset15_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg335_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg336_in = par_reset15_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg336_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg337_in = par_reset15_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg337_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg338_in = par_reset15_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg338_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_done_reg339_in = par_reset15_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd15 & !par_reset15_out & go) ? 1'd1 : '0;
  assign par_done_reg339_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd15 & !par_reset15_out & go | par_reset15_out) ? 1'd1 : '0;
  assign par_reset16_in = par_reset16_out ? 1'd0 : (par_done_reg340_out & par_done_reg341_out & par_done_reg342_out & par_done_reg343_out & par_done_reg344_out & par_done_reg345_out & par_done_reg346_out & par_done_reg347_out & par_done_reg348_out & par_done_reg349_out & par_done_reg350_out & par_done_reg351_out & par_done_reg352_out & par_done_reg353_out & par_done_reg354_out & par_done_reg355_out & par_done_reg356_out & par_done_reg357_out & par_done_reg358_out & par_done_reg359_out & par_done_reg360_out & par_done_reg361_out & par_done_reg362_out & par_done_reg363_out & par_done_reg364_out & par_done_reg365_out & par_done_reg366_out & par_done_reg367_out & par_done_reg368_out & par_done_reg369_out & par_done_reg370_out & par_done_reg371_out & par_done_reg372_out & par_done_reg373_out & par_done_reg374_out & par_done_reg375_out & par_done_reg376_out & par_done_reg377_out & par_done_reg378_out & par_done_reg379_out & par_done_reg380_out & par_done_reg381_out & par_done_reg382_out & par_done_reg383_out & par_done_reg384_out & par_done_reg385_out & par_done_reg386_out & par_done_reg387_out & par_done_reg388_out & par_done_reg389_out & par_done_reg390_out & par_done_reg391_out & par_done_reg392_out & par_done_reg393_out & par_done_reg394_out & par_done_reg395_out & par_done_reg396_out & par_done_reg397_out & par_done_reg398_out & par_done_reg399_out & par_done_reg400_out & par_done_reg401_out & par_done_reg402_out & par_done_reg403_out & par_done_reg404_out & par_done_reg405_out & par_done_reg406_out & par_done_reg407_out & par_done_reg408_out & par_done_reg409_out & par_done_reg410_out & par_done_reg411_out & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_reset16_write_en = (par_done_reg340_out & par_done_reg341_out & par_done_reg342_out & par_done_reg343_out & par_done_reg344_out & par_done_reg345_out & par_done_reg346_out & par_done_reg347_out & par_done_reg348_out & par_done_reg349_out & par_done_reg350_out & par_done_reg351_out & par_done_reg352_out & par_done_reg353_out & par_done_reg354_out & par_done_reg355_out & par_done_reg356_out & par_done_reg357_out & par_done_reg358_out & par_done_reg359_out & par_done_reg360_out & par_done_reg361_out & par_done_reg362_out & par_done_reg363_out & par_done_reg364_out & par_done_reg365_out & par_done_reg366_out & par_done_reg367_out & par_done_reg368_out & par_done_reg369_out & par_done_reg370_out & par_done_reg371_out & par_done_reg372_out & par_done_reg373_out & par_done_reg374_out & par_done_reg375_out & par_done_reg376_out & par_done_reg377_out & par_done_reg378_out & par_done_reg379_out & par_done_reg380_out & par_done_reg381_out & par_done_reg382_out & par_done_reg383_out & par_done_reg384_out & par_done_reg385_out & par_done_reg386_out & par_done_reg387_out & par_done_reg388_out & par_done_reg389_out & par_done_reg390_out & par_done_reg391_out & par_done_reg392_out & par_done_reg393_out & par_done_reg394_out & par_done_reg395_out & par_done_reg396_out & par_done_reg397_out & par_done_reg398_out & par_done_reg399_out & par_done_reg400_out & par_done_reg401_out & par_done_reg402_out & par_done_reg403_out & par_done_reg404_out & par_done_reg405_out & par_done_reg406_out & par_done_reg407_out & par_done_reg408_out & par_done_reg409_out & par_done_reg410_out & par_done_reg411_out & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg340_in = par_reset16_out ? 1'd0 : (top_00_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg340_write_en = (top_00_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg341_in = par_reset16_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg341_write_en = (top_01_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg342_in = par_reset16_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg342_write_en = (top_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg343_in = par_reset16_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg343_write_en = (top_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg344_in = par_reset16_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg344_write_en = (top_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg345_in = par_reset16_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg345_write_en = (top_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg346_in = par_reset16_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg346_write_en = (top_06_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg347_in = par_reset16_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg347_write_en = (top_07_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg348_in = par_reset16_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg348_write_en = (top_10_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg349_in = par_reset16_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg349_write_en = (top_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg350_in = par_reset16_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg350_write_en = (top_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg351_in = par_reset16_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg351_write_en = (top_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg352_in = par_reset16_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg352_write_en = (top_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg353_in = par_reset16_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg353_write_en = (top_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg354_in = par_reset16_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg354_write_en = (top_16_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg355_in = par_reset16_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg355_write_en = (top_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg356_in = par_reset16_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg356_write_en = (top_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg357_in = par_reset16_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg357_write_en = (top_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg358_in = par_reset16_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg358_write_en = (top_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg359_in = par_reset16_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg359_write_en = (top_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg360_in = par_reset16_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg360_write_en = (top_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg361_in = par_reset16_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg361_write_en = (top_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg362_in = par_reset16_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg362_write_en = (top_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg363_in = par_reset16_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg363_write_en = (top_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg364_in = par_reset16_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg364_write_en = (top_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg365_in = par_reset16_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg365_write_en = (top_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg366_in = par_reset16_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg366_write_en = (top_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg367_in = par_reset16_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg367_write_en = (top_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg368_in = par_reset16_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg368_write_en = (top_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg369_in = par_reset16_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg369_write_en = (top_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg370_in = par_reset16_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg370_write_en = (top_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg371_in = par_reset16_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg371_write_en = (top_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg372_in = par_reset16_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg372_write_en = (top_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg373_in = par_reset16_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg373_write_en = (top_60_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg374_in = par_reset16_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg374_write_en = (top_61_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg375_in = par_reset16_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg375_write_en = (top_70_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg376_in = par_reset16_out ? 1'd0 : (left_00_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg376_write_en = (left_00_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg377_in = par_reset16_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg377_write_en = (left_01_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg378_in = par_reset16_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg378_write_en = (left_02_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg379_in = par_reset16_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg379_write_en = (left_03_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg380_in = par_reset16_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg380_write_en = (left_04_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg381_in = par_reset16_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg381_write_en = (left_05_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg382_in = par_reset16_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg382_write_en = (left_06_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg383_in = par_reset16_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg383_write_en = (left_07_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg384_in = par_reset16_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg384_write_en = (left_10_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg385_in = par_reset16_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg385_write_en = (left_11_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg386_in = par_reset16_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg386_write_en = (left_12_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg387_in = par_reset16_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg387_write_en = (left_13_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg388_in = par_reset16_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg388_write_en = (left_14_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg389_in = par_reset16_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg389_write_en = (left_15_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg390_in = par_reset16_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg390_write_en = (left_16_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg391_in = par_reset16_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg391_write_en = (left_20_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg392_in = par_reset16_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg392_write_en = (left_21_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg393_in = par_reset16_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg393_write_en = (left_22_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg394_in = par_reset16_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg394_write_en = (left_23_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg395_in = par_reset16_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg395_write_en = (left_24_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg396_in = par_reset16_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg396_write_en = (left_25_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg397_in = par_reset16_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg397_write_en = (left_30_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg398_in = par_reset16_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg398_write_en = (left_31_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg399_in = par_reset16_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg399_write_en = (left_32_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg400_in = par_reset16_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg400_write_en = (left_33_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg401_in = par_reset16_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg401_write_en = (left_34_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg402_in = par_reset16_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg402_write_en = (left_40_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg403_in = par_reset16_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg403_write_en = (left_41_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg404_in = par_reset16_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg404_write_en = (left_42_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg405_in = par_reset16_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg405_write_en = (left_43_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg406_in = par_reset16_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg406_write_en = (left_50_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg407_in = par_reset16_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg407_write_en = (left_51_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg408_in = par_reset16_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg408_write_en = (left_52_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg409_in = par_reset16_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg409_write_en = (left_60_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg410_in = par_reset16_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg410_write_en = (left_61_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_done_reg411_in = par_reset16_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd16 & !par_reset16_out & go) ? 1'd1 : '0;
  assign par_done_reg411_write_en = (left_70_read_done & fsm0_out == 32'd16 & !par_reset16_out & go | par_reset16_out) ? 1'd1 : '0;
  assign par_reset17_in = par_reset17_out ? 1'd0 : (par_done_reg412_out & par_done_reg413_out & par_done_reg414_out & par_done_reg415_out & par_done_reg416_out & par_done_reg417_out & par_done_reg418_out & par_done_reg419_out & par_done_reg420_out & par_done_reg421_out & par_done_reg422_out & par_done_reg423_out & par_done_reg424_out & par_done_reg425_out & par_done_reg426_out & par_done_reg427_out & par_done_reg428_out & par_done_reg429_out & par_done_reg430_out & par_done_reg431_out & par_done_reg432_out & par_done_reg433_out & par_done_reg434_out & par_done_reg435_out & par_done_reg436_out & par_done_reg437_out & par_done_reg438_out & par_done_reg439_out & par_done_reg440_out & par_done_reg441_out & par_done_reg442_out & par_done_reg443_out & par_done_reg444_out & par_done_reg445_out & par_done_reg446_out & par_done_reg447_out & par_done_reg448_out & par_done_reg449_out & par_done_reg450_out & par_done_reg451_out & par_done_reg452_out & par_done_reg453_out & par_done_reg454_out & par_done_reg455_out & par_done_reg456_out & par_done_reg457_out & par_done_reg458_out & par_done_reg459_out & par_done_reg460_out & par_done_reg461_out & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_reset17_write_en = (par_done_reg412_out & par_done_reg413_out & par_done_reg414_out & par_done_reg415_out & par_done_reg416_out & par_done_reg417_out & par_done_reg418_out & par_done_reg419_out & par_done_reg420_out & par_done_reg421_out & par_done_reg422_out & par_done_reg423_out & par_done_reg424_out & par_done_reg425_out & par_done_reg426_out & par_done_reg427_out & par_done_reg428_out & par_done_reg429_out & par_done_reg430_out & par_done_reg431_out & par_done_reg432_out & par_done_reg433_out & par_done_reg434_out & par_done_reg435_out & par_done_reg436_out & par_done_reg437_out & par_done_reg438_out & par_done_reg439_out & par_done_reg440_out & par_done_reg441_out & par_done_reg442_out & par_done_reg443_out & par_done_reg444_out & par_done_reg445_out & par_done_reg446_out & par_done_reg447_out & par_done_reg448_out & par_done_reg449_out & par_done_reg450_out & par_done_reg451_out & par_done_reg452_out & par_done_reg453_out & par_done_reg454_out & par_done_reg455_out & par_done_reg456_out & par_done_reg457_out & par_done_reg458_out & par_done_reg459_out & par_done_reg460_out & par_done_reg461_out & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg412_in = par_reset17_out ? 1'd0 : (t1_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg412_write_en = (t1_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg413_in = par_reset17_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg413_write_en = (t2_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg414_in = par_reset17_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg414_write_en = (t3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg415_in = par_reset17_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg415_write_en = (t4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg416_in = par_reset17_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg416_write_en = (t5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg417_in = par_reset17_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg417_write_en = (t6_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg418_in = par_reset17_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg418_write_en = (t7_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg419_in = par_reset17_out ? 1'd0 : (l1_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg419_write_en = (l1_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg420_in = par_reset17_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg420_write_en = (l2_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg421_in = par_reset17_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg421_write_en = (l3_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg422_in = par_reset17_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg422_write_en = (l4_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg423_in = par_reset17_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg423_write_en = (l5_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg424_in = par_reset17_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg424_write_en = (l6_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg425_in = par_reset17_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg425_write_en = (l7_idx_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg426_in = par_reset17_out ? 1'd0 : (right_00_write_done & down_00_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg426_write_en = (right_00_write_done & down_00_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg427_in = par_reset17_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg427_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg428_in = par_reset17_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg428_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg429_in = par_reset17_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg429_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg430_in = par_reset17_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg430_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg431_in = par_reset17_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg431_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg432_in = par_reset17_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg432_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg433_in = par_reset17_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg433_write_en = (down_07_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg434_in = par_reset17_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg434_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg435_in = par_reset17_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg435_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg436_in = par_reset17_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg436_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg437_in = par_reset17_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg437_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg438_in = par_reset17_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg438_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg439_in = par_reset17_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg439_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg440_in = par_reset17_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg440_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg441_in = par_reset17_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg441_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg442_in = par_reset17_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg442_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg443_in = par_reset17_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg443_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg444_in = par_reset17_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg444_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg445_in = par_reset17_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg445_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg446_in = par_reset17_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg446_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg447_in = par_reset17_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg447_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg448_in = par_reset17_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg448_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg449_in = par_reset17_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg449_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg450_in = par_reset17_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg450_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg451_in = par_reset17_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg451_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg452_in = par_reset17_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg452_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg453_in = par_reset17_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg453_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg454_in = par_reset17_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg454_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg455_in = par_reset17_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg455_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg456_in = par_reset17_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg456_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg457_in = par_reset17_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg457_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg458_in = par_reset17_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg458_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg459_in = par_reset17_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg459_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg460_in = par_reset17_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg460_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_done_reg461_in = par_reset17_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd17 & !par_reset17_out & go) ? 1'd1 : '0;
  assign par_done_reg461_write_en = (right_70_write_done & fsm0_out == 32'd17 & !par_reset17_out & go | par_reset17_out) ? 1'd1 : '0;
  assign par_reset18_in = par_reset18_out ? 1'd0 : (par_done_reg462_out & par_done_reg463_out & par_done_reg464_out & par_done_reg465_out & par_done_reg466_out & par_done_reg467_out & par_done_reg468_out & par_done_reg469_out & par_done_reg470_out & par_done_reg471_out & par_done_reg472_out & par_done_reg473_out & par_done_reg474_out & par_done_reg475_out & par_done_reg476_out & par_done_reg477_out & par_done_reg478_out & par_done_reg479_out & par_done_reg480_out & par_done_reg481_out & par_done_reg482_out & par_done_reg483_out & par_done_reg484_out & par_done_reg485_out & par_done_reg486_out & par_done_reg487_out & par_done_reg488_out & par_done_reg489_out & par_done_reg490_out & par_done_reg491_out & par_done_reg492_out & par_done_reg493_out & par_done_reg494_out & par_done_reg495_out & par_done_reg496_out & par_done_reg497_out & par_done_reg498_out & par_done_reg499_out & par_done_reg500_out & par_done_reg501_out & par_done_reg502_out & par_done_reg503_out & par_done_reg504_out & par_done_reg505_out & par_done_reg506_out & par_done_reg507_out & par_done_reg508_out & par_done_reg509_out & par_done_reg510_out & par_done_reg511_out & par_done_reg512_out & par_done_reg513_out & par_done_reg514_out & par_done_reg515_out & par_done_reg516_out & par_done_reg517_out & par_done_reg518_out & par_done_reg519_out & par_done_reg520_out & par_done_reg521_out & par_done_reg522_out & par_done_reg523_out & par_done_reg524_out & par_done_reg525_out & par_done_reg526_out & par_done_reg527_out & par_done_reg528_out & par_done_reg529_out & par_done_reg530_out & par_done_reg531_out & par_done_reg532_out & par_done_reg533_out & par_done_reg534_out & par_done_reg535_out & par_done_reg536_out & par_done_reg537_out & par_done_reg538_out & par_done_reg539_out & par_done_reg540_out & par_done_reg541_out & par_done_reg542_out & par_done_reg543_out & par_done_reg544_out & par_done_reg545_out & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_reset18_write_en = (par_done_reg462_out & par_done_reg463_out & par_done_reg464_out & par_done_reg465_out & par_done_reg466_out & par_done_reg467_out & par_done_reg468_out & par_done_reg469_out & par_done_reg470_out & par_done_reg471_out & par_done_reg472_out & par_done_reg473_out & par_done_reg474_out & par_done_reg475_out & par_done_reg476_out & par_done_reg477_out & par_done_reg478_out & par_done_reg479_out & par_done_reg480_out & par_done_reg481_out & par_done_reg482_out & par_done_reg483_out & par_done_reg484_out & par_done_reg485_out & par_done_reg486_out & par_done_reg487_out & par_done_reg488_out & par_done_reg489_out & par_done_reg490_out & par_done_reg491_out & par_done_reg492_out & par_done_reg493_out & par_done_reg494_out & par_done_reg495_out & par_done_reg496_out & par_done_reg497_out & par_done_reg498_out & par_done_reg499_out & par_done_reg500_out & par_done_reg501_out & par_done_reg502_out & par_done_reg503_out & par_done_reg504_out & par_done_reg505_out & par_done_reg506_out & par_done_reg507_out & par_done_reg508_out & par_done_reg509_out & par_done_reg510_out & par_done_reg511_out & par_done_reg512_out & par_done_reg513_out & par_done_reg514_out & par_done_reg515_out & par_done_reg516_out & par_done_reg517_out & par_done_reg518_out & par_done_reg519_out & par_done_reg520_out & par_done_reg521_out & par_done_reg522_out & par_done_reg523_out & par_done_reg524_out & par_done_reg525_out & par_done_reg526_out & par_done_reg527_out & par_done_reg528_out & par_done_reg529_out & par_done_reg530_out & par_done_reg531_out & par_done_reg532_out & par_done_reg533_out & par_done_reg534_out & par_done_reg535_out & par_done_reg536_out & par_done_reg537_out & par_done_reg538_out & par_done_reg539_out & par_done_reg540_out & par_done_reg541_out & par_done_reg542_out & par_done_reg543_out & par_done_reg544_out & par_done_reg545_out & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg462_in = par_reset18_out ? 1'd0 : (top_01_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg462_write_en = (top_01_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg463_in = par_reset18_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg463_write_en = (top_02_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg464_in = par_reset18_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg464_write_en = (top_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg465_in = par_reset18_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg465_write_en = (top_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg466_in = par_reset18_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg466_write_en = (top_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg467_in = par_reset18_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg467_write_en = (top_06_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg468_in = par_reset18_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg468_write_en = (top_07_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg469_in = par_reset18_out ? 1'd0 : (top_10_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg469_write_en = (top_10_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg470_in = par_reset18_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg470_write_en = (top_11_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg471_in = par_reset18_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg471_write_en = (top_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg472_in = par_reset18_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg472_write_en = (top_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg473_in = par_reset18_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg473_write_en = (top_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg474_in = par_reset18_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg474_write_en = (top_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg475_in = par_reset18_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg475_write_en = (top_16_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg476_in = par_reset18_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg476_write_en = (top_17_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg477_in = par_reset18_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg477_write_en = (top_20_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg478_in = par_reset18_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg478_write_en = (top_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg479_in = par_reset18_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg479_write_en = (top_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg480_in = par_reset18_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg480_write_en = (top_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg481_in = par_reset18_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg481_write_en = (top_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg482_in = par_reset18_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg482_write_en = (top_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg483_in = par_reset18_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg483_write_en = (top_26_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg484_in = par_reset18_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg484_write_en = (top_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg485_in = par_reset18_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg485_write_en = (top_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg486_in = par_reset18_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg486_write_en = (top_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg487_in = par_reset18_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg487_write_en = (top_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg488_in = par_reset18_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg488_write_en = (top_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg489_in = par_reset18_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg489_write_en = (top_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg490_in = par_reset18_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg490_write_en = (top_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg491_in = par_reset18_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg491_write_en = (top_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg492_in = par_reset18_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg492_write_en = (top_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg493_in = par_reset18_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg493_write_en = (top_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg494_in = par_reset18_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg494_write_en = (top_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg495_in = par_reset18_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg495_write_en = (top_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg496_in = par_reset18_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg496_write_en = (top_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg497_in = par_reset18_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg497_write_en = (top_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg498_in = par_reset18_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg498_write_en = (top_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg499_in = par_reset18_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg499_write_en = (top_60_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg500_in = par_reset18_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg500_write_en = (top_61_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg501_in = par_reset18_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg501_write_en = (top_62_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg502_in = par_reset18_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg502_write_en = (top_70_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg503_in = par_reset18_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg503_write_en = (top_71_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg504_in = par_reset18_out ? 1'd0 : (left_01_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg504_write_en = (left_01_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg505_in = par_reset18_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg505_write_en = (left_02_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg506_in = par_reset18_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg506_write_en = (left_03_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg507_in = par_reset18_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg507_write_en = (left_04_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg508_in = par_reset18_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg508_write_en = (left_05_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg509_in = par_reset18_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg509_write_en = (left_06_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg510_in = par_reset18_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg510_write_en = (left_07_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg511_in = par_reset18_out ? 1'd0 : (left_10_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg511_write_en = (left_10_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg512_in = par_reset18_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg512_write_en = (left_11_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg513_in = par_reset18_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg513_write_en = (left_12_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg514_in = par_reset18_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg514_write_en = (left_13_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg515_in = par_reset18_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg515_write_en = (left_14_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg516_in = par_reset18_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg516_write_en = (left_15_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg517_in = par_reset18_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg517_write_en = (left_16_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg518_in = par_reset18_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg518_write_en = (left_17_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg519_in = par_reset18_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg519_write_en = (left_20_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg520_in = par_reset18_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg520_write_en = (left_21_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg521_in = par_reset18_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg521_write_en = (left_22_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg522_in = par_reset18_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg522_write_en = (left_23_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg523_in = par_reset18_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg523_write_en = (left_24_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg524_in = par_reset18_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg524_write_en = (left_25_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg525_in = par_reset18_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg525_write_en = (left_26_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg526_in = par_reset18_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg526_write_en = (left_30_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg527_in = par_reset18_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg527_write_en = (left_31_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg528_in = par_reset18_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg528_write_en = (left_32_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg529_in = par_reset18_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg529_write_en = (left_33_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg530_in = par_reset18_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg530_write_en = (left_34_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg531_in = par_reset18_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg531_write_en = (left_35_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg532_in = par_reset18_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg532_write_en = (left_40_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg533_in = par_reset18_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg533_write_en = (left_41_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg534_in = par_reset18_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg534_write_en = (left_42_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg535_in = par_reset18_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg535_write_en = (left_43_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg536_in = par_reset18_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg536_write_en = (left_44_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg537_in = par_reset18_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg537_write_en = (left_50_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg538_in = par_reset18_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg538_write_en = (left_51_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg539_in = par_reset18_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg539_write_en = (left_52_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg540_in = par_reset18_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg540_write_en = (left_53_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg541_in = par_reset18_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg541_write_en = (left_60_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg542_in = par_reset18_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg542_write_en = (left_61_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg543_in = par_reset18_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg543_write_en = (left_62_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg544_in = par_reset18_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg544_write_en = (left_70_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_done_reg545_in = par_reset18_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd18 & !par_reset18_out & go) ? 1'd1 : '0;
  assign par_done_reg545_write_en = (left_71_read_done & fsm0_out == 32'd18 & !par_reset18_out & go | par_reset18_out) ? 1'd1 : '0;
  assign par_reset19_in = par_reset19_out ? 1'd0 : (par_done_reg546_out & par_done_reg547_out & par_done_reg548_out & par_done_reg549_out & par_done_reg550_out & par_done_reg551_out & par_done_reg552_out & par_done_reg553_out & par_done_reg554_out & par_done_reg555_out & par_done_reg556_out & par_done_reg557_out & par_done_reg558_out & par_done_reg559_out & par_done_reg560_out & par_done_reg561_out & par_done_reg562_out & par_done_reg563_out & par_done_reg564_out & par_done_reg565_out & par_done_reg566_out & par_done_reg567_out & par_done_reg568_out & par_done_reg569_out & par_done_reg570_out & par_done_reg571_out & par_done_reg572_out & par_done_reg573_out & par_done_reg574_out & par_done_reg575_out & par_done_reg576_out & par_done_reg577_out & par_done_reg578_out & par_done_reg579_out & par_done_reg580_out & par_done_reg581_out & par_done_reg582_out & par_done_reg583_out & par_done_reg584_out & par_done_reg585_out & par_done_reg586_out & par_done_reg587_out & par_done_reg588_out & par_done_reg589_out & par_done_reg590_out & par_done_reg591_out & par_done_reg592_out & par_done_reg593_out & par_done_reg594_out & par_done_reg595_out & par_done_reg596_out & par_done_reg597_out & par_done_reg598_out & par_done_reg599_out & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_reset19_write_en = (par_done_reg546_out & par_done_reg547_out & par_done_reg548_out & par_done_reg549_out & par_done_reg550_out & par_done_reg551_out & par_done_reg552_out & par_done_reg553_out & par_done_reg554_out & par_done_reg555_out & par_done_reg556_out & par_done_reg557_out & par_done_reg558_out & par_done_reg559_out & par_done_reg560_out & par_done_reg561_out & par_done_reg562_out & par_done_reg563_out & par_done_reg564_out & par_done_reg565_out & par_done_reg566_out & par_done_reg567_out & par_done_reg568_out & par_done_reg569_out & par_done_reg570_out & par_done_reg571_out & par_done_reg572_out & par_done_reg573_out & par_done_reg574_out & par_done_reg575_out & par_done_reg576_out & par_done_reg577_out & par_done_reg578_out & par_done_reg579_out & par_done_reg580_out & par_done_reg581_out & par_done_reg582_out & par_done_reg583_out & par_done_reg584_out & par_done_reg585_out & par_done_reg586_out & par_done_reg587_out & par_done_reg588_out & par_done_reg589_out & par_done_reg590_out & par_done_reg591_out & par_done_reg592_out & par_done_reg593_out & par_done_reg594_out & par_done_reg595_out & par_done_reg596_out & par_done_reg597_out & par_done_reg598_out & par_done_reg599_out & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg546_in = par_reset19_out ? 1'd0 : (t2_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg546_write_en = (t2_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg547_in = par_reset19_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg547_write_en = (t3_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg548_in = par_reset19_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg548_write_en = (t4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg549_in = par_reset19_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg549_write_en = (t5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg550_in = par_reset19_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg550_write_en = (t6_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg551_in = par_reset19_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg551_write_en = (t7_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg552_in = par_reset19_out ? 1'd0 : (l2_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg552_write_en = (l2_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg553_in = par_reset19_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg553_write_en = (l3_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg554_in = par_reset19_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg554_write_en = (l4_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg555_in = par_reset19_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg555_write_en = (l5_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg556_in = par_reset19_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg556_write_en = (l6_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg557_in = par_reset19_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg557_write_en = (l7_idx_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg558_in = par_reset19_out ? 1'd0 : (right_01_write_done & down_01_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg558_write_en = (right_01_write_done & down_01_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg559_in = par_reset19_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg559_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg560_in = par_reset19_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg560_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg561_in = par_reset19_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg561_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg562_in = par_reset19_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg562_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg563_in = par_reset19_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg563_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg564_in = par_reset19_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg564_write_en = (down_07_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg565_in = par_reset19_out ? 1'd0 : (right_10_write_done & down_10_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg565_write_en = (right_10_write_done & down_10_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg566_in = par_reset19_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg566_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg567_in = par_reset19_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg567_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg568_in = par_reset19_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg568_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg569_in = par_reset19_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg569_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg570_in = par_reset19_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg570_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg571_in = par_reset19_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg571_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg572_in = par_reset19_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg572_write_en = (down_17_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg573_in = par_reset19_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg573_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg574_in = par_reset19_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg574_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg575_in = par_reset19_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg575_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg576_in = par_reset19_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg576_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg577_in = par_reset19_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg577_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg578_in = par_reset19_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg578_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg579_in = par_reset19_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg579_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg580_in = par_reset19_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg580_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg581_in = par_reset19_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg581_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg582_in = par_reset19_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg582_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg583_in = par_reset19_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg583_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg584_in = par_reset19_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg584_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg585_in = par_reset19_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg585_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg586_in = par_reset19_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg586_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg587_in = par_reset19_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg587_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg588_in = par_reset19_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg588_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg589_in = par_reset19_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg589_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg590_in = par_reset19_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg590_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg591_in = par_reset19_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg591_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg592_in = par_reset19_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg592_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg593_in = par_reset19_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg593_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg594_in = par_reset19_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg594_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg595_in = par_reset19_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg595_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg596_in = par_reset19_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg596_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg597_in = par_reset19_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg597_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg598_in = par_reset19_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg598_write_en = (right_70_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_done_reg599_in = par_reset19_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd19 & !par_reset19_out & go) ? 1'd1 : '0;
  assign par_done_reg599_write_en = (right_71_write_done & fsm0_out == 32'd19 & !par_reset19_out & go | par_reset19_out) ? 1'd1 : '0;
  assign par_reset20_in = par_reset20_out ? 1'd0 : (par_done_reg600_out & par_done_reg601_out & par_done_reg602_out & par_done_reg603_out & par_done_reg604_out & par_done_reg605_out & par_done_reg606_out & par_done_reg607_out & par_done_reg608_out & par_done_reg609_out & par_done_reg610_out & par_done_reg611_out & par_done_reg612_out & par_done_reg613_out & par_done_reg614_out & par_done_reg615_out & par_done_reg616_out & par_done_reg617_out & par_done_reg618_out & par_done_reg619_out & par_done_reg620_out & par_done_reg621_out & par_done_reg622_out & par_done_reg623_out & par_done_reg624_out & par_done_reg625_out & par_done_reg626_out & par_done_reg627_out & par_done_reg628_out & par_done_reg629_out & par_done_reg630_out & par_done_reg631_out & par_done_reg632_out & par_done_reg633_out & par_done_reg634_out & par_done_reg635_out & par_done_reg636_out & par_done_reg637_out & par_done_reg638_out & par_done_reg639_out & par_done_reg640_out & par_done_reg641_out & par_done_reg642_out & par_done_reg643_out & par_done_reg644_out & par_done_reg645_out & par_done_reg646_out & par_done_reg647_out & par_done_reg648_out & par_done_reg649_out & par_done_reg650_out & par_done_reg651_out & par_done_reg652_out & par_done_reg653_out & par_done_reg654_out & par_done_reg655_out & par_done_reg656_out & par_done_reg657_out & par_done_reg658_out & par_done_reg659_out & par_done_reg660_out & par_done_reg661_out & par_done_reg662_out & par_done_reg663_out & par_done_reg664_out & par_done_reg665_out & par_done_reg666_out & par_done_reg667_out & par_done_reg668_out & par_done_reg669_out & par_done_reg670_out & par_done_reg671_out & par_done_reg672_out & par_done_reg673_out & par_done_reg674_out & par_done_reg675_out & par_done_reg676_out & par_done_reg677_out & par_done_reg678_out & par_done_reg679_out & par_done_reg680_out & par_done_reg681_out & par_done_reg682_out & par_done_reg683_out & par_done_reg684_out & par_done_reg685_out & par_done_reg686_out & par_done_reg687_out & par_done_reg688_out & par_done_reg689_out & par_done_reg690_out & par_done_reg691_out & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_reset20_write_en = (par_done_reg600_out & par_done_reg601_out & par_done_reg602_out & par_done_reg603_out & par_done_reg604_out & par_done_reg605_out & par_done_reg606_out & par_done_reg607_out & par_done_reg608_out & par_done_reg609_out & par_done_reg610_out & par_done_reg611_out & par_done_reg612_out & par_done_reg613_out & par_done_reg614_out & par_done_reg615_out & par_done_reg616_out & par_done_reg617_out & par_done_reg618_out & par_done_reg619_out & par_done_reg620_out & par_done_reg621_out & par_done_reg622_out & par_done_reg623_out & par_done_reg624_out & par_done_reg625_out & par_done_reg626_out & par_done_reg627_out & par_done_reg628_out & par_done_reg629_out & par_done_reg630_out & par_done_reg631_out & par_done_reg632_out & par_done_reg633_out & par_done_reg634_out & par_done_reg635_out & par_done_reg636_out & par_done_reg637_out & par_done_reg638_out & par_done_reg639_out & par_done_reg640_out & par_done_reg641_out & par_done_reg642_out & par_done_reg643_out & par_done_reg644_out & par_done_reg645_out & par_done_reg646_out & par_done_reg647_out & par_done_reg648_out & par_done_reg649_out & par_done_reg650_out & par_done_reg651_out & par_done_reg652_out & par_done_reg653_out & par_done_reg654_out & par_done_reg655_out & par_done_reg656_out & par_done_reg657_out & par_done_reg658_out & par_done_reg659_out & par_done_reg660_out & par_done_reg661_out & par_done_reg662_out & par_done_reg663_out & par_done_reg664_out & par_done_reg665_out & par_done_reg666_out & par_done_reg667_out & par_done_reg668_out & par_done_reg669_out & par_done_reg670_out & par_done_reg671_out & par_done_reg672_out & par_done_reg673_out & par_done_reg674_out & par_done_reg675_out & par_done_reg676_out & par_done_reg677_out & par_done_reg678_out & par_done_reg679_out & par_done_reg680_out & par_done_reg681_out & par_done_reg682_out & par_done_reg683_out & par_done_reg684_out & par_done_reg685_out & par_done_reg686_out & par_done_reg687_out & par_done_reg688_out & par_done_reg689_out & par_done_reg690_out & par_done_reg691_out & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg600_in = par_reset20_out ? 1'd0 : (top_02_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg600_write_en = (top_02_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg601_in = par_reset20_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg601_write_en = (top_03_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg602_in = par_reset20_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg602_write_en = (top_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg603_in = par_reset20_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg603_write_en = (top_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg604_in = par_reset20_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg604_write_en = (top_06_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg605_in = par_reset20_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg605_write_en = (top_07_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg606_in = par_reset20_out ? 1'd0 : (top_11_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg606_write_en = (top_11_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg607_in = par_reset20_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg607_write_en = (top_12_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg608_in = par_reset20_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg608_write_en = (top_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg609_in = par_reset20_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg609_write_en = (top_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg610_in = par_reset20_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg610_write_en = (top_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg611_in = par_reset20_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg611_write_en = (top_16_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg612_in = par_reset20_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg612_write_en = (top_17_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg613_in = par_reset20_out ? 1'd0 : (top_20_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg613_write_en = (top_20_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg614_in = par_reset20_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg614_write_en = (top_21_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg615_in = par_reset20_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg615_write_en = (top_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg616_in = par_reset20_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg616_write_en = (top_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg617_in = par_reset20_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg617_write_en = (top_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg618_in = par_reset20_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg618_write_en = (top_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg619_in = par_reset20_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg619_write_en = (top_26_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg620_in = par_reset20_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg620_write_en = (top_27_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg621_in = par_reset20_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg621_write_en = (top_30_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg622_in = par_reset20_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg622_write_en = (top_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg623_in = par_reset20_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg623_write_en = (top_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg624_in = par_reset20_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg624_write_en = (top_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg625_in = par_reset20_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg625_write_en = (top_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg626_in = par_reset20_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg626_write_en = (top_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg627_in = par_reset20_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg627_write_en = (top_36_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg628_in = par_reset20_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg628_write_en = (top_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg629_in = par_reset20_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg629_write_en = (top_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg630_in = par_reset20_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg630_write_en = (top_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg631_in = par_reset20_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg631_write_en = (top_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg632_in = par_reset20_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg632_write_en = (top_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg633_in = par_reset20_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg633_write_en = (top_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg634_in = par_reset20_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg634_write_en = (top_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg635_in = par_reset20_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg635_write_en = (top_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg636_in = par_reset20_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg636_write_en = (top_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg637_in = par_reset20_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg637_write_en = (top_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg638_in = par_reset20_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg638_write_en = (top_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg639_in = par_reset20_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg639_write_en = (top_60_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg640_in = par_reset20_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg640_write_en = (top_61_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg641_in = par_reset20_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg641_write_en = (top_62_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg642_in = par_reset20_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg642_write_en = (top_63_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg643_in = par_reset20_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg643_write_en = (top_70_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg644_in = par_reset20_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg644_write_en = (top_71_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg645_in = par_reset20_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg645_write_en = (top_72_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg646_in = par_reset20_out ? 1'd0 : (left_02_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg646_write_en = (left_02_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg647_in = par_reset20_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg647_write_en = (left_03_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg648_in = par_reset20_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg648_write_en = (left_04_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg649_in = par_reset20_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg649_write_en = (left_05_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg650_in = par_reset20_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg650_write_en = (left_06_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg651_in = par_reset20_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg651_write_en = (left_07_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg652_in = par_reset20_out ? 1'd0 : (left_11_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg652_write_en = (left_11_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg653_in = par_reset20_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg653_write_en = (left_12_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg654_in = par_reset20_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg654_write_en = (left_13_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg655_in = par_reset20_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg655_write_en = (left_14_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg656_in = par_reset20_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg656_write_en = (left_15_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg657_in = par_reset20_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg657_write_en = (left_16_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg658_in = par_reset20_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg658_write_en = (left_17_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg659_in = par_reset20_out ? 1'd0 : (left_20_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg659_write_en = (left_20_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg660_in = par_reset20_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg660_write_en = (left_21_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg661_in = par_reset20_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg661_write_en = (left_22_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg662_in = par_reset20_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg662_write_en = (left_23_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg663_in = par_reset20_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg663_write_en = (left_24_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg664_in = par_reset20_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg664_write_en = (left_25_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg665_in = par_reset20_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg665_write_en = (left_26_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg666_in = par_reset20_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg666_write_en = (left_27_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg667_in = par_reset20_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg667_write_en = (left_30_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg668_in = par_reset20_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg668_write_en = (left_31_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg669_in = par_reset20_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg669_write_en = (left_32_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg670_in = par_reset20_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg670_write_en = (left_33_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg671_in = par_reset20_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg671_write_en = (left_34_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg672_in = par_reset20_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg672_write_en = (left_35_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg673_in = par_reset20_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg673_write_en = (left_36_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg674_in = par_reset20_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg674_write_en = (left_40_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg675_in = par_reset20_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg675_write_en = (left_41_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg676_in = par_reset20_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg676_write_en = (left_42_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg677_in = par_reset20_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg677_write_en = (left_43_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg678_in = par_reset20_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg678_write_en = (left_44_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg679_in = par_reset20_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg679_write_en = (left_45_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg680_in = par_reset20_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg680_write_en = (left_50_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg681_in = par_reset20_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg681_write_en = (left_51_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg682_in = par_reset20_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg682_write_en = (left_52_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg683_in = par_reset20_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg683_write_en = (left_53_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg684_in = par_reset20_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg684_write_en = (left_54_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg685_in = par_reset20_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg685_write_en = (left_60_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg686_in = par_reset20_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg686_write_en = (left_61_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg687_in = par_reset20_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg687_write_en = (left_62_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg688_in = par_reset20_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg688_write_en = (left_63_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg689_in = par_reset20_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg689_write_en = (left_70_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg690_in = par_reset20_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg690_write_en = (left_71_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_done_reg691_in = par_reset20_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd20 & !par_reset20_out & go) ? 1'd1 : '0;
  assign par_done_reg691_write_en = (left_72_read_done & fsm0_out == 32'd20 & !par_reset20_out & go | par_reset20_out) ? 1'd1 : '0;
  assign par_reset21_in = par_reset21_out ? 1'd0 : (par_done_reg692_out & par_done_reg693_out & par_done_reg694_out & par_done_reg695_out & par_done_reg696_out & par_done_reg697_out & par_done_reg698_out & par_done_reg699_out & par_done_reg700_out & par_done_reg701_out & par_done_reg702_out & par_done_reg703_out & par_done_reg704_out & par_done_reg705_out & par_done_reg706_out & par_done_reg707_out & par_done_reg708_out & par_done_reg709_out & par_done_reg710_out & par_done_reg711_out & par_done_reg712_out & par_done_reg713_out & par_done_reg714_out & par_done_reg715_out & par_done_reg716_out & par_done_reg717_out & par_done_reg718_out & par_done_reg719_out & par_done_reg720_out & par_done_reg721_out & par_done_reg722_out & par_done_reg723_out & par_done_reg724_out & par_done_reg725_out & par_done_reg726_out & par_done_reg727_out & par_done_reg728_out & par_done_reg729_out & par_done_reg730_out & par_done_reg731_out & par_done_reg732_out & par_done_reg733_out & par_done_reg734_out & par_done_reg735_out & par_done_reg736_out & par_done_reg737_out & par_done_reg738_out & par_done_reg739_out & par_done_reg740_out & par_done_reg741_out & par_done_reg742_out & par_done_reg743_out & par_done_reg744_out & par_done_reg745_out & par_done_reg746_out & par_done_reg747_out & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_reset21_write_en = (par_done_reg692_out & par_done_reg693_out & par_done_reg694_out & par_done_reg695_out & par_done_reg696_out & par_done_reg697_out & par_done_reg698_out & par_done_reg699_out & par_done_reg700_out & par_done_reg701_out & par_done_reg702_out & par_done_reg703_out & par_done_reg704_out & par_done_reg705_out & par_done_reg706_out & par_done_reg707_out & par_done_reg708_out & par_done_reg709_out & par_done_reg710_out & par_done_reg711_out & par_done_reg712_out & par_done_reg713_out & par_done_reg714_out & par_done_reg715_out & par_done_reg716_out & par_done_reg717_out & par_done_reg718_out & par_done_reg719_out & par_done_reg720_out & par_done_reg721_out & par_done_reg722_out & par_done_reg723_out & par_done_reg724_out & par_done_reg725_out & par_done_reg726_out & par_done_reg727_out & par_done_reg728_out & par_done_reg729_out & par_done_reg730_out & par_done_reg731_out & par_done_reg732_out & par_done_reg733_out & par_done_reg734_out & par_done_reg735_out & par_done_reg736_out & par_done_reg737_out & par_done_reg738_out & par_done_reg739_out & par_done_reg740_out & par_done_reg741_out & par_done_reg742_out & par_done_reg743_out & par_done_reg744_out & par_done_reg745_out & par_done_reg746_out & par_done_reg747_out & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg692_in = par_reset21_out ? 1'd0 : (t3_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg692_write_en = (t3_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg693_in = par_reset21_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg693_write_en = (t4_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg694_in = par_reset21_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg694_write_en = (t5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg695_in = par_reset21_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg695_write_en = (t6_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg696_in = par_reset21_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg696_write_en = (t7_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg697_in = par_reset21_out ? 1'd0 : (l3_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg697_write_en = (l3_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg698_in = par_reset21_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg698_write_en = (l4_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg699_in = par_reset21_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg699_write_en = (l5_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg700_in = par_reset21_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg700_write_en = (l6_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg701_in = par_reset21_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg701_write_en = (l7_idx_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg702_in = par_reset21_out ? 1'd0 : (right_02_write_done & down_02_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg702_write_en = (right_02_write_done & down_02_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg703_in = par_reset21_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg703_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg704_in = par_reset21_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg704_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg705_in = par_reset21_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg705_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg706_in = par_reset21_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg706_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg707_in = par_reset21_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg707_write_en = (down_07_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg708_in = par_reset21_out ? 1'd0 : (right_11_write_done & down_11_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg708_write_en = (right_11_write_done & down_11_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg709_in = par_reset21_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg709_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg710_in = par_reset21_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg710_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg711_in = par_reset21_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg711_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg712_in = par_reset21_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg712_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg713_in = par_reset21_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg713_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg714_in = par_reset21_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg714_write_en = (down_17_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg715_in = par_reset21_out ? 1'd0 : (right_20_write_done & down_20_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg715_write_en = (right_20_write_done & down_20_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg716_in = par_reset21_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg716_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg717_in = par_reset21_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg717_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg718_in = par_reset21_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg718_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg719_in = par_reset21_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg719_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg720_in = par_reset21_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg720_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg721_in = par_reset21_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg721_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg722_in = par_reset21_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg722_write_en = (down_27_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg723_in = par_reset21_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg723_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg724_in = par_reset21_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg724_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg725_in = par_reset21_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg725_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg726_in = par_reset21_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg726_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg727_in = par_reset21_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg727_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg728_in = par_reset21_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg728_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg729_in = par_reset21_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg729_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg730_in = par_reset21_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg730_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg731_in = par_reset21_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg731_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg732_in = par_reset21_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg732_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg733_in = par_reset21_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg733_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg734_in = par_reset21_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg734_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg735_in = par_reset21_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg735_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg736_in = par_reset21_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg736_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg737_in = par_reset21_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg737_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg738_in = par_reset21_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg738_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg739_in = par_reset21_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg739_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg740_in = par_reset21_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg740_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg741_in = par_reset21_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg741_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg742_in = par_reset21_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg742_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg743_in = par_reset21_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg743_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg744_in = par_reset21_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg744_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg745_in = par_reset21_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg745_write_en = (right_70_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg746_in = par_reset21_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg746_write_en = (right_71_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_done_reg747_in = par_reset21_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd21 & !par_reset21_out & go) ? 1'd1 : '0;
  assign par_done_reg747_write_en = (right_72_write_done & fsm0_out == 32'd21 & !par_reset21_out & go | par_reset21_out) ? 1'd1 : '0;
  assign par_reset22_in = par_reset22_out ? 1'd0 : (par_done_reg748_out & par_done_reg749_out & par_done_reg750_out & par_done_reg751_out & par_done_reg752_out & par_done_reg753_out & par_done_reg754_out & par_done_reg755_out & par_done_reg756_out & par_done_reg757_out & par_done_reg758_out & par_done_reg759_out & par_done_reg760_out & par_done_reg761_out & par_done_reg762_out & par_done_reg763_out & par_done_reg764_out & par_done_reg765_out & par_done_reg766_out & par_done_reg767_out & par_done_reg768_out & par_done_reg769_out & par_done_reg770_out & par_done_reg771_out & par_done_reg772_out & par_done_reg773_out & par_done_reg774_out & par_done_reg775_out & par_done_reg776_out & par_done_reg777_out & par_done_reg778_out & par_done_reg779_out & par_done_reg780_out & par_done_reg781_out & par_done_reg782_out & par_done_reg783_out & par_done_reg784_out & par_done_reg785_out & par_done_reg786_out & par_done_reg787_out & par_done_reg788_out & par_done_reg789_out & par_done_reg790_out & par_done_reg791_out & par_done_reg792_out & par_done_reg793_out & par_done_reg794_out & par_done_reg795_out & par_done_reg796_out & par_done_reg797_out & par_done_reg798_out & par_done_reg799_out & par_done_reg800_out & par_done_reg801_out & par_done_reg802_out & par_done_reg803_out & par_done_reg804_out & par_done_reg805_out & par_done_reg806_out & par_done_reg807_out & par_done_reg808_out & par_done_reg809_out & par_done_reg810_out & par_done_reg811_out & par_done_reg812_out & par_done_reg813_out & par_done_reg814_out & par_done_reg815_out & par_done_reg816_out & par_done_reg817_out & par_done_reg818_out & par_done_reg819_out & par_done_reg820_out & par_done_reg821_out & par_done_reg822_out & par_done_reg823_out & par_done_reg824_out & par_done_reg825_out & par_done_reg826_out & par_done_reg827_out & par_done_reg828_out & par_done_reg829_out & par_done_reg830_out & par_done_reg831_out & par_done_reg832_out & par_done_reg833_out & par_done_reg834_out & par_done_reg835_out & par_done_reg836_out & par_done_reg837_out & par_done_reg838_out & par_done_reg839_out & par_done_reg840_out & par_done_reg841_out & par_done_reg842_out & par_done_reg843_out & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_reset22_write_en = (par_done_reg748_out & par_done_reg749_out & par_done_reg750_out & par_done_reg751_out & par_done_reg752_out & par_done_reg753_out & par_done_reg754_out & par_done_reg755_out & par_done_reg756_out & par_done_reg757_out & par_done_reg758_out & par_done_reg759_out & par_done_reg760_out & par_done_reg761_out & par_done_reg762_out & par_done_reg763_out & par_done_reg764_out & par_done_reg765_out & par_done_reg766_out & par_done_reg767_out & par_done_reg768_out & par_done_reg769_out & par_done_reg770_out & par_done_reg771_out & par_done_reg772_out & par_done_reg773_out & par_done_reg774_out & par_done_reg775_out & par_done_reg776_out & par_done_reg777_out & par_done_reg778_out & par_done_reg779_out & par_done_reg780_out & par_done_reg781_out & par_done_reg782_out & par_done_reg783_out & par_done_reg784_out & par_done_reg785_out & par_done_reg786_out & par_done_reg787_out & par_done_reg788_out & par_done_reg789_out & par_done_reg790_out & par_done_reg791_out & par_done_reg792_out & par_done_reg793_out & par_done_reg794_out & par_done_reg795_out & par_done_reg796_out & par_done_reg797_out & par_done_reg798_out & par_done_reg799_out & par_done_reg800_out & par_done_reg801_out & par_done_reg802_out & par_done_reg803_out & par_done_reg804_out & par_done_reg805_out & par_done_reg806_out & par_done_reg807_out & par_done_reg808_out & par_done_reg809_out & par_done_reg810_out & par_done_reg811_out & par_done_reg812_out & par_done_reg813_out & par_done_reg814_out & par_done_reg815_out & par_done_reg816_out & par_done_reg817_out & par_done_reg818_out & par_done_reg819_out & par_done_reg820_out & par_done_reg821_out & par_done_reg822_out & par_done_reg823_out & par_done_reg824_out & par_done_reg825_out & par_done_reg826_out & par_done_reg827_out & par_done_reg828_out & par_done_reg829_out & par_done_reg830_out & par_done_reg831_out & par_done_reg832_out & par_done_reg833_out & par_done_reg834_out & par_done_reg835_out & par_done_reg836_out & par_done_reg837_out & par_done_reg838_out & par_done_reg839_out & par_done_reg840_out & par_done_reg841_out & par_done_reg842_out & par_done_reg843_out & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg748_in = par_reset22_out ? 1'd0 : (top_03_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg748_write_en = (top_03_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg749_in = par_reset22_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg749_write_en = (top_04_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg750_in = par_reset22_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg750_write_en = (top_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg751_in = par_reset22_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg751_write_en = (top_06_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg752_in = par_reset22_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg752_write_en = (top_07_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg753_in = par_reset22_out ? 1'd0 : (top_12_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg753_write_en = (top_12_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg754_in = par_reset22_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg754_write_en = (top_13_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg755_in = par_reset22_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg755_write_en = (top_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg756_in = par_reset22_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg756_write_en = (top_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg757_in = par_reset22_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg757_write_en = (top_16_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg758_in = par_reset22_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg758_write_en = (top_17_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg759_in = par_reset22_out ? 1'd0 : (top_21_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg759_write_en = (top_21_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg760_in = par_reset22_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg760_write_en = (top_22_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg761_in = par_reset22_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg761_write_en = (top_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg762_in = par_reset22_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg762_write_en = (top_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg763_in = par_reset22_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg763_write_en = (top_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg764_in = par_reset22_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg764_write_en = (top_26_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg765_in = par_reset22_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg765_write_en = (top_27_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg766_in = par_reset22_out ? 1'd0 : (top_30_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg766_write_en = (top_30_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg767_in = par_reset22_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg767_write_en = (top_31_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg768_in = par_reset22_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg768_write_en = (top_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg769_in = par_reset22_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg769_write_en = (top_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg770_in = par_reset22_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg770_write_en = (top_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg771_in = par_reset22_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg771_write_en = (top_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg772_in = par_reset22_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg772_write_en = (top_36_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg773_in = par_reset22_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg773_write_en = (top_37_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg774_in = par_reset22_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg774_write_en = (top_40_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg775_in = par_reset22_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg775_write_en = (top_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg776_in = par_reset22_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg776_write_en = (top_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg777_in = par_reset22_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg777_write_en = (top_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg778_in = par_reset22_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg778_write_en = (top_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg779_in = par_reset22_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg779_write_en = (top_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg780_in = par_reset22_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg780_write_en = (top_46_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg781_in = par_reset22_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg781_write_en = (top_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg782_in = par_reset22_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg782_write_en = (top_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg783_in = par_reset22_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg783_write_en = (top_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg784_in = par_reset22_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg784_write_en = (top_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg785_in = par_reset22_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg785_write_en = (top_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg786_in = par_reset22_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg786_write_en = (top_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg787_in = par_reset22_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg787_write_en = (top_60_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg788_in = par_reset22_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg788_write_en = (top_61_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg789_in = par_reset22_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg789_write_en = (top_62_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg790_in = par_reset22_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg790_write_en = (top_63_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg791_in = par_reset22_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg791_write_en = (top_64_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg792_in = par_reset22_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg792_write_en = (top_70_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg793_in = par_reset22_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg793_write_en = (top_71_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg794_in = par_reset22_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg794_write_en = (top_72_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg795_in = par_reset22_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg795_write_en = (top_73_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg796_in = par_reset22_out ? 1'd0 : (left_03_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg796_write_en = (left_03_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg797_in = par_reset22_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg797_write_en = (left_04_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg798_in = par_reset22_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg798_write_en = (left_05_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg799_in = par_reset22_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg799_write_en = (left_06_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg800_in = par_reset22_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg800_write_en = (left_07_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg801_in = par_reset22_out ? 1'd0 : (left_12_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg801_write_en = (left_12_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg802_in = par_reset22_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg802_write_en = (left_13_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg803_in = par_reset22_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg803_write_en = (left_14_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg804_in = par_reset22_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg804_write_en = (left_15_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg805_in = par_reset22_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg805_write_en = (left_16_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg806_in = par_reset22_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg806_write_en = (left_17_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg807_in = par_reset22_out ? 1'd0 : (left_21_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg807_write_en = (left_21_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg808_in = par_reset22_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg808_write_en = (left_22_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg809_in = par_reset22_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg809_write_en = (left_23_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg810_in = par_reset22_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg810_write_en = (left_24_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg811_in = par_reset22_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg811_write_en = (left_25_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg812_in = par_reset22_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg812_write_en = (left_26_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg813_in = par_reset22_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg813_write_en = (left_27_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg814_in = par_reset22_out ? 1'd0 : (left_30_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg814_write_en = (left_30_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg815_in = par_reset22_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg815_write_en = (left_31_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg816_in = par_reset22_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg816_write_en = (left_32_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg817_in = par_reset22_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg817_write_en = (left_33_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg818_in = par_reset22_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg818_write_en = (left_34_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg819_in = par_reset22_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg819_write_en = (left_35_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg820_in = par_reset22_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg820_write_en = (left_36_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg821_in = par_reset22_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg821_write_en = (left_37_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg822_in = par_reset22_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg822_write_en = (left_40_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg823_in = par_reset22_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg823_write_en = (left_41_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg824_in = par_reset22_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg824_write_en = (left_42_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg825_in = par_reset22_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg825_write_en = (left_43_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg826_in = par_reset22_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg826_write_en = (left_44_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg827_in = par_reset22_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg827_write_en = (left_45_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg828_in = par_reset22_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg828_write_en = (left_46_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg829_in = par_reset22_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg829_write_en = (left_50_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg830_in = par_reset22_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg830_write_en = (left_51_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg831_in = par_reset22_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg831_write_en = (left_52_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg832_in = par_reset22_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg832_write_en = (left_53_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg833_in = par_reset22_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg833_write_en = (left_54_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg834_in = par_reset22_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg834_write_en = (left_55_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg835_in = par_reset22_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg835_write_en = (left_60_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg836_in = par_reset22_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg836_write_en = (left_61_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg837_in = par_reset22_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg837_write_en = (left_62_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg838_in = par_reset22_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg838_write_en = (left_63_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg839_in = par_reset22_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg839_write_en = (left_64_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg840_in = par_reset22_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg840_write_en = (left_70_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg841_in = par_reset22_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg841_write_en = (left_71_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg842_in = par_reset22_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg842_write_en = (left_72_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_done_reg843_in = par_reset22_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd22 & !par_reset22_out & go) ? 1'd1 : '0;
  assign par_done_reg843_write_en = (left_73_read_done & fsm0_out == 32'd22 & !par_reset22_out & go | par_reset22_out) ? 1'd1 : '0;
  assign par_reset23_in = par_reset23_out ? 1'd0 : (par_done_reg844_out & par_done_reg845_out & par_done_reg846_out & par_done_reg847_out & par_done_reg848_out & par_done_reg849_out & par_done_reg850_out & par_done_reg851_out & par_done_reg852_out & par_done_reg853_out & par_done_reg854_out & par_done_reg855_out & par_done_reg856_out & par_done_reg857_out & par_done_reg858_out & par_done_reg859_out & par_done_reg860_out & par_done_reg861_out & par_done_reg862_out & par_done_reg863_out & par_done_reg864_out & par_done_reg865_out & par_done_reg866_out & par_done_reg867_out & par_done_reg868_out & par_done_reg869_out & par_done_reg870_out & par_done_reg871_out & par_done_reg872_out & par_done_reg873_out & par_done_reg874_out & par_done_reg875_out & par_done_reg876_out & par_done_reg877_out & par_done_reg878_out & par_done_reg879_out & par_done_reg880_out & par_done_reg881_out & par_done_reg882_out & par_done_reg883_out & par_done_reg884_out & par_done_reg885_out & par_done_reg886_out & par_done_reg887_out & par_done_reg888_out & par_done_reg889_out & par_done_reg890_out & par_done_reg891_out & par_done_reg892_out & par_done_reg893_out & par_done_reg894_out & par_done_reg895_out & par_done_reg896_out & par_done_reg897_out & par_done_reg898_out & par_done_reg899_out & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_reset23_write_en = (par_done_reg844_out & par_done_reg845_out & par_done_reg846_out & par_done_reg847_out & par_done_reg848_out & par_done_reg849_out & par_done_reg850_out & par_done_reg851_out & par_done_reg852_out & par_done_reg853_out & par_done_reg854_out & par_done_reg855_out & par_done_reg856_out & par_done_reg857_out & par_done_reg858_out & par_done_reg859_out & par_done_reg860_out & par_done_reg861_out & par_done_reg862_out & par_done_reg863_out & par_done_reg864_out & par_done_reg865_out & par_done_reg866_out & par_done_reg867_out & par_done_reg868_out & par_done_reg869_out & par_done_reg870_out & par_done_reg871_out & par_done_reg872_out & par_done_reg873_out & par_done_reg874_out & par_done_reg875_out & par_done_reg876_out & par_done_reg877_out & par_done_reg878_out & par_done_reg879_out & par_done_reg880_out & par_done_reg881_out & par_done_reg882_out & par_done_reg883_out & par_done_reg884_out & par_done_reg885_out & par_done_reg886_out & par_done_reg887_out & par_done_reg888_out & par_done_reg889_out & par_done_reg890_out & par_done_reg891_out & par_done_reg892_out & par_done_reg893_out & par_done_reg894_out & par_done_reg895_out & par_done_reg896_out & par_done_reg897_out & par_done_reg898_out & par_done_reg899_out & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg844_in = par_reset23_out ? 1'd0 : (t4_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg844_write_en = (t4_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg845_in = par_reset23_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg845_write_en = (t5_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg846_in = par_reset23_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg846_write_en = (t6_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg847_in = par_reset23_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg847_write_en = (t7_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg848_in = par_reset23_out ? 1'd0 : (l4_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg848_write_en = (l4_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg849_in = par_reset23_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg849_write_en = (l5_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg850_in = par_reset23_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg850_write_en = (l6_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg851_in = par_reset23_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg851_write_en = (l7_idx_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg852_in = par_reset23_out ? 1'd0 : (right_03_write_done & down_03_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg852_write_en = (right_03_write_done & down_03_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg853_in = par_reset23_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg853_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg854_in = par_reset23_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg854_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg855_in = par_reset23_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg855_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg856_in = par_reset23_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg856_write_en = (down_07_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg857_in = par_reset23_out ? 1'd0 : (right_12_write_done & down_12_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg857_write_en = (right_12_write_done & down_12_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg858_in = par_reset23_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg858_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg859_in = par_reset23_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg859_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg860_in = par_reset23_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg860_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg861_in = par_reset23_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg861_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg862_in = par_reset23_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg862_write_en = (down_17_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg863_in = par_reset23_out ? 1'd0 : (right_21_write_done & down_21_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg863_write_en = (right_21_write_done & down_21_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg864_in = par_reset23_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg864_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg865_in = par_reset23_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg865_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg866_in = par_reset23_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg866_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg867_in = par_reset23_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg867_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg868_in = par_reset23_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg868_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg869_in = par_reset23_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg869_write_en = (down_27_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg870_in = par_reset23_out ? 1'd0 : (right_30_write_done & down_30_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg870_write_en = (right_30_write_done & down_30_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg871_in = par_reset23_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg871_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg872_in = par_reset23_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg872_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg873_in = par_reset23_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg873_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg874_in = par_reset23_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg874_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg875_in = par_reset23_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg875_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg876_in = par_reset23_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg876_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg877_in = par_reset23_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg877_write_en = (down_37_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg878_in = par_reset23_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg878_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg879_in = par_reset23_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg879_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg880_in = par_reset23_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg880_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg881_in = par_reset23_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg881_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg882_in = par_reset23_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg882_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg883_in = par_reset23_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg883_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg884_in = par_reset23_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg884_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg885_in = par_reset23_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg885_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg886_in = par_reset23_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg886_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg887_in = par_reset23_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg887_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg888_in = par_reset23_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg888_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg889_in = par_reset23_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg889_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg890_in = par_reset23_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg890_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg891_in = par_reset23_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg891_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg892_in = par_reset23_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg892_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg893_in = par_reset23_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg893_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg894_in = par_reset23_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg894_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg895_in = par_reset23_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg895_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg896_in = par_reset23_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg896_write_en = (right_70_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg897_in = par_reset23_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg897_write_en = (right_71_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg898_in = par_reset23_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg898_write_en = (right_72_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_done_reg899_in = par_reset23_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd23 & !par_reset23_out & go) ? 1'd1 : '0;
  assign par_done_reg899_write_en = (right_73_write_done & fsm0_out == 32'd23 & !par_reset23_out & go | par_reset23_out) ? 1'd1 : '0;
  assign par_reset24_in = par_reset24_out ? 1'd0 : (par_done_reg900_out & par_done_reg901_out & par_done_reg902_out & par_done_reg903_out & par_done_reg904_out & par_done_reg905_out & par_done_reg906_out & par_done_reg907_out & par_done_reg908_out & par_done_reg909_out & par_done_reg910_out & par_done_reg911_out & par_done_reg912_out & par_done_reg913_out & par_done_reg914_out & par_done_reg915_out & par_done_reg916_out & par_done_reg917_out & par_done_reg918_out & par_done_reg919_out & par_done_reg920_out & par_done_reg921_out & par_done_reg922_out & par_done_reg923_out & par_done_reg924_out & par_done_reg925_out & par_done_reg926_out & par_done_reg927_out & par_done_reg928_out & par_done_reg929_out & par_done_reg930_out & par_done_reg931_out & par_done_reg932_out & par_done_reg933_out & par_done_reg934_out & par_done_reg935_out & par_done_reg936_out & par_done_reg937_out & par_done_reg938_out & par_done_reg939_out & par_done_reg940_out & par_done_reg941_out & par_done_reg942_out & par_done_reg943_out & par_done_reg944_out & par_done_reg945_out & par_done_reg946_out & par_done_reg947_out & par_done_reg948_out & par_done_reg949_out & par_done_reg950_out & par_done_reg951_out & par_done_reg952_out & par_done_reg953_out & par_done_reg954_out & par_done_reg955_out & par_done_reg956_out & par_done_reg957_out & par_done_reg958_out & par_done_reg959_out & par_done_reg960_out & par_done_reg961_out & par_done_reg962_out & par_done_reg963_out & par_done_reg964_out & par_done_reg965_out & par_done_reg966_out & par_done_reg967_out & par_done_reg968_out & par_done_reg969_out & par_done_reg970_out & par_done_reg971_out & par_done_reg972_out & par_done_reg973_out & par_done_reg974_out & par_done_reg975_out & par_done_reg976_out & par_done_reg977_out & par_done_reg978_out & par_done_reg979_out & par_done_reg980_out & par_done_reg981_out & par_done_reg982_out & par_done_reg983_out & par_done_reg984_out & par_done_reg985_out & par_done_reg986_out & par_done_reg987_out & par_done_reg988_out & par_done_reg989_out & par_done_reg990_out & par_done_reg991_out & par_done_reg992_out & par_done_reg993_out & par_done_reg994_out & par_done_reg995_out & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_reset24_write_en = (par_done_reg900_out & par_done_reg901_out & par_done_reg902_out & par_done_reg903_out & par_done_reg904_out & par_done_reg905_out & par_done_reg906_out & par_done_reg907_out & par_done_reg908_out & par_done_reg909_out & par_done_reg910_out & par_done_reg911_out & par_done_reg912_out & par_done_reg913_out & par_done_reg914_out & par_done_reg915_out & par_done_reg916_out & par_done_reg917_out & par_done_reg918_out & par_done_reg919_out & par_done_reg920_out & par_done_reg921_out & par_done_reg922_out & par_done_reg923_out & par_done_reg924_out & par_done_reg925_out & par_done_reg926_out & par_done_reg927_out & par_done_reg928_out & par_done_reg929_out & par_done_reg930_out & par_done_reg931_out & par_done_reg932_out & par_done_reg933_out & par_done_reg934_out & par_done_reg935_out & par_done_reg936_out & par_done_reg937_out & par_done_reg938_out & par_done_reg939_out & par_done_reg940_out & par_done_reg941_out & par_done_reg942_out & par_done_reg943_out & par_done_reg944_out & par_done_reg945_out & par_done_reg946_out & par_done_reg947_out & par_done_reg948_out & par_done_reg949_out & par_done_reg950_out & par_done_reg951_out & par_done_reg952_out & par_done_reg953_out & par_done_reg954_out & par_done_reg955_out & par_done_reg956_out & par_done_reg957_out & par_done_reg958_out & par_done_reg959_out & par_done_reg960_out & par_done_reg961_out & par_done_reg962_out & par_done_reg963_out & par_done_reg964_out & par_done_reg965_out & par_done_reg966_out & par_done_reg967_out & par_done_reg968_out & par_done_reg969_out & par_done_reg970_out & par_done_reg971_out & par_done_reg972_out & par_done_reg973_out & par_done_reg974_out & par_done_reg975_out & par_done_reg976_out & par_done_reg977_out & par_done_reg978_out & par_done_reg979_out & par_done_reg980_out & par_done_reg981_out & par_done_reg982_out & par_done_reg983_out & par_done_reg984_out & par_done_reg985_out & par_done_reg986_out & par_done_reg987_out & par_done_reg988_out & par_done_reg989_out & par_done_reg990_out & par_done_reg991_out & par_done_reg992_out & par_done_reg993_out & par_done_reg994_out & par_done_reg995_out & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg900_in = par_reset24_out ? 1'd0 : (top_04_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg900_write_en = (top_04_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg901_in = par_reset24_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg901_write_en = (top_05_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg902_in = par_reset24_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg902_write_en = (top_06_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg903_in = par_reset24_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg903_write_en = (top_07_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg904_in = par_reset24_out ? 1'd0 : (top_13_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg904_write_en = (top_13_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg905_in = par_reset24_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg905_write_en = (top_14_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg906_in = par_reset24_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg906_write_en = (top_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg907_in = par_reset24_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg907_write_en = (top_16_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg908_in = par_reset24_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg908_write_en = (top_17_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg909_in = par_reset24_out ? 1'd0 : (top_22_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg909_write_en = (top_22_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg910_in = par_reset24_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg910_write_en = (top_23_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg911_in = par_reset24_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg911_write_en = (top_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg912_in = par_reset24_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg912_write_en = (top_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg913_in = par_reset24_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg913_write_en = (top_26_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg914_in = par_reset24_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg914_write_en = (top_27_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg915_in = par_reset24_out ? 1'd0 : (top_31_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg915_write_en = (top_31_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg916_in = par_reset24_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg916_write_en = (top_32_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg917_in = par_reset24_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg917_write_en = (top_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg918_in = par_reset24_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg918_write_en = (top_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg919_in = par_reset24_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg919_write_en = (top_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg920_in = par_reset24_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg920_write_en = (top_36_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg921_in = par_reset24_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg921_write_en = (top_37_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg922_in = par_reset24_out ? 1'd0 : (top_40_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg922_write_en = (top_40_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg923_in = par_reset24_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg923_write_en = (top_41_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg924_in = par_reset24_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg924_write_en = (top_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg925_in = par_reset24_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg925_write_en = (top_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg926_in = par_reset24_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg926_write_en = (top_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg927_in = par_reset24_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg927_write_en = (top_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg928_in = par_reset24_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg928_write_en = (top_46_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg929_in = par_reset24_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg929_write_en = (top_47_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg930_in = par_reset24_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg930_write_en = (top_50_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg931_in = par_reset24_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg931_write_en = (top_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg932_in = par_reset24_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg932_write_en = (top_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg933_in = par_reset24_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg933_write_en = (top_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg934_in = par_reset24_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg934_write_en = (top_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg935_in = par_reset24_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg935_write_en = (top_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg936_in = par_reset24_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg936_write_en = (top_56_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg937_in = par_reset24_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg937_write_en = (top_60_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg938_in = par_reset24_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg938_write_en = (top_61_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg939_in = par_reset24_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg939_write_en = (top_62_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg940_in = par_reset24_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg940_write_en = (top_63_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg941_in = par_reset24_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg941_write_en = (top_64_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg942_in = par_reset24_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg942_write_en = (top_65_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg943_in = par_reset24_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg943_write_en = (top_70_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg944_in = par_reset24_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg944_write_en = (top_71_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg945_in = par_reset24_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg945_write_en = (top_72_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg946_in = par_reset24_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg946_write_en = (top_73_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg947_in = par_reset24_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg947_write_en = (top_74_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg948_in = par_reset24_out ? 1'd0 : (left_04_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg948_write_en = (left_04_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg949_in = par_reset24_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg949_write_en = (left_05_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg950_in = par_reset24_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg950_write_en = (left_06_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg951_in = par_reset24_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg951_write_en = (left_07_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg952_in = par_reset24_out ? 1'd0 : (left_13_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg952_write_en = (left_13_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg953_in = par_reset24_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg953_write_en = (left_14_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg954_in = par_reset24_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg954_write_en = (left_15_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg955_in = par_reset24_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg955_write_en = (left_16_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg956_in = par_reset24_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg956_write_en = (left_17_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg957_in = par_reset24_out ? 1'd0 : (left_22_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg957_write_en = (left_22_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg958_in = par_reset24_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg958_write_en = (left_23_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg959_in = par_reset24_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg959_write_en = (left_24_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg960_in = par_reset24_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg960_write_en = (left_25_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg961_in = par_reset24_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg961_write_en = (left_26_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg962_in = par_reset24_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg962_write_en = (left_27_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg963_in = par_reset24_out ? 1'd0 : (left_31_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg963_write_en = (left_31_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg964_in = par_reset24_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg964_write_en = (left_32_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg965_in = par_reset24_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg965_write_en = (left_33_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg966_in = par_reset24_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg966_write_en = (left_34_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg967_in = par_reset24_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg967_write_en = (left_35_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg968_in = par_reset24_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg968_write_en = (left_36_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg969_in = par_reset24_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg969_write_en = (left_37_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg970_in = par_reset24_out ? 1'd0 : (left_40_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg970_write_en = (left_40_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg971_in = par_reset24_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg971_write_en = (left_41_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg972_in = par_reset24_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg972_write_en = (left_42_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg973_in = par_reset24_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg973_write_en = (left_43_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg974_in = par_reset24_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg974_write_en = (left_44_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg975_in = par_reset24_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg975_write_en = (left_45_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg976_in = par_reset24_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg976_write_en = (left_46_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg977_in = par_reset24_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg977_write_en = (left_47_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg978_in = par_reset24_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg978_write_en = (left_50_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg979_in = par_reset24_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg979_write_en = (left_51_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg980_in = par_reset24_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg980_write_en = (left_52_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg981_in = par_reset24_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg981_write_en = (left_53_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg982_in = par_reset24_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg982_write_en = (left_54_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg983_in = par_reset24_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg983_write_en = (left_55_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg984_in = par_reset24_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg984_write_en = (left_56_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg985_in = par_reset24_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg985_write_en = (left_60_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg986_in = par_reset24_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg986_write_en = (left_61_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg987_in = par_reset24_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg987_write_en = (left_62_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg988_in = par_reset24_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg988_write_en = (left_63_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg989_in = par_reset24_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg989_write_en = (left_64_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg990_in = par_reset24_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg990_write_en = (left_65_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg991_in = par_reset24_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg991_write_en = (left_70_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg992_in = par_reset24_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg992_write_en = (left_71_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg993_in = par_reset24_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg993_write_en = (left_72_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg994_in = par_reset24_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg994_write_en = (left_73_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_done_reg995_in = par_reset24_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd24 & !par_reset24_out & go) ? 1'd1 : '0;
  assign par_done_reg995_write_en = (left_74_read_done & fsm0_out == 32'd24 & !par_reset24_out & go | par_reset24_out) ? 1'd1 : '0;
  assign par_reset25_in = par_reset25_out ? 1'd0 : (par_done_reg996_out & par_done_reg997_out & par_done_reg998_out & par_done_reg999_out & par_done_reg1000_out & par_done_reg1001_out & par_done_reg1002_out & par_done_reg1003_out & par_done_reg1004_out & par_done_reg1005_out & par_done_reg1006_out & par_done_reg1007_out & par_done_reg1008_out & par_done_reg1009_out & par_done_reg1010_out & par_done_reg1011_out & par_done_reg1012_out & par_done_reg1013_out & par_done_reg1014_out & par_done_reg1015_out & par_done_reg1016_out & par_done_reg1017_out & par_done_reg1018_out & par_done_reg1019_out & par_done_reg1020_out & par_done_reg1021_out & par_done_reg1022_out & par_done_reg1023_out & par_done_reg1024_out & par_done_reg1025_out & par_done_reg1026_out & par_done_reg1027_out & par_done_reg1028_out & par_done_reg1029_out & par_done_reg1030_out & par_done_reg1031_out & par_done_reg1032_out & par_done_reg1033_out & par_done_reg1034_out & par_done_reg1035_out & par_done_reg1036_out & par_done_reg1037_out & par_done_reg1038_out & par_done_reg1039_out & par_done_reg1040_out & par_done_reg1041_out & par_done_reg1042_out & par_done_reg1043_out & par_done_reg1044_out & par_done_reg1045_out & par_done_reg1046_out & par_done_reg1047_out & par_done_reg1048_out & par_done_reg1049_out & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_reset25_write_en = (par_done_reg996_out & par_done_reg997_out & par_done_reg998_out & par_done_reg999_out & par_done_reg1000_out & par_done_reg1001_out & par_done_reg1002_out & par_done_reg1003_out & par_done_reg1004_out & par_done_reg1005_out & par_done_reg1006_out & par_done_reg1007_out & par_done_reg1008_out & par_done_reg1009_out & par_done_reg1010_out & par_done_reg1011_out & par_done_reg1012_out & par_done_reg1013_out & par_done_reg1014_out & par_done_reg1015_out & par_done_reg1016_out & par_done_reg1017_out & par_done_reg1018_out & par_done_reg1019_out & par_done_reg1020_out & par_done_reg1021_out & par_done_reg1022_out & par_done_reg1023_out & par_done_reg1024_out & par_done_reg1025_out & par_done_reg1026_out & par_done_reg1027_out & par_done_reg1028_out & par_done_reg1029_out & par_done_reg1030_out & par_done_reg1031_out & par_done_reg1032_out & par_done_reg1033_out & par_done_reg1034_out & par_done_reg1035_out & par_done_reg1036_out & par_done_reg1037_out & par_done_reg1038_out & par_done_reg1039_out & par_done_reg1040_out & par_done_reg1041_out & par_done_reg1042_out & par_done_reg1043_out & par_done_reg1044_out & par_done_reg1045_out & par_done_reg1046_out & par_done_reg1047_out & par_done_reg1048_out & par_done_reg1049_out & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg996_in = par_reset25_out ? 1'd0 : (t5_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg996_write_en = (t5_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg997_in = par_reset25_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg997_write_en = (t6_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg998_in = par_reset25_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg998_write_en = (t7_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg999_in = par_reset25_out ? 1'd0 : (l5_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg999_write_en = (l5_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1000_in = par_reset25_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1000_write_en = (l6_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1001_in = par_reset25_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1001_write_en = (l7_idx_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1002_in = par_reset25_out ? 1'd0 : (right_04_write_done & down_04_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1002_write_en = (right_04_write_done & down_04_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1003_in = par_reset25_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1003_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1004_in = par_reset25_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1004_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1005_in = par_reset25_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1005_write_en = (down_07_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1006_in = par_reset25_out ? 1'd0 : (right_13_write_done & down_13_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1006_write_en = (right_13_write_done & down_13_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1007_in = par_reset25_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1007_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1008_in = par_reset25_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1008_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1009_in = par_reset25_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1009_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1010_in = par_reset25_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1010_write_en = (down_17_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1011_in = par_reset25_out ? 1'd0 : (right_22_write_done & down_22_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1011_write_en = (right_22_write_done & down_22_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1012_in = par_reset25_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1012_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1013_in = par_reset25_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1013_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1014_in = par_reset25_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1014_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1015_in = par_reset25_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1015_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1016_in = par_reset25_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1016_write_en = (down_27_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1017_in = par_reset25_out ? 1'd0 : (right_31_write_done & down_31_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1017_write_en = (right_31_write_done & down_31_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1018_in = par_reset25_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1018_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1019_in = par_reset25_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1019_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1020_in = par_reset25_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1020_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1021_in = par_reset25_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1021_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1022_in = par_reset25_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1022_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1023_in = par_reset25_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1023_write_en = (down_37_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1024_in = par_reset25_out ? 1'd0 : (right_40_write_done & down_40_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1024_write_en = (right_40_write_done & down_40_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1025_in = par_reset25_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1025_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1026_in = par_reset25_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1026_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1027_in = par_reset25_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1027_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1028_in = par_reset25_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1028_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1029_in = par_reset25_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1029_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1030_in = par_reset25_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1030_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1031_in = par_reset25_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1031_write_en = (down_47_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1032_in = par_reset25_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1032_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1033_in = par_reset25_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1033_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1034_in = par_reset25_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1034_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1035_in = par_reset25_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1035_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1036_in = par_reset25_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1036_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1037_in = par_reset25_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1037_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1038_in = par_reset25_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1038_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1039_in = par_reset25_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1039_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1040_in = par_reset25_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1040_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1041_in = par_reset25_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1041_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1042_in = par_reset25_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1042_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1043_in = par_reset25_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1043_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1044_in = par_reset25_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1044_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1045_in = par_reset25_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1045_write_en = (right_70_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1046_in = par_reset25_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1046_write_en = (right_71_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1047_in = par_reset25_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1047_write_en = (right_72_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1048_in = par_reset25_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1048_write_en = (right_73_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_done_reg1049_in = par_reset25_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd25 & !par_reset25_out & go) ? 1'd1 : '0;
  assign par_done_reg1049_write_en = (right_74_write_done & fsm0_out == 32'd25 & !par_reset25_out & go | par_reset25_out) ? 1'd1 : '0;
  assign par_reset26_in = par_reset26_out ? 1'd0 : (par_done_reg1050_out & par_done_reg1051_out & par_done_reg1052_out & par_done_reg1053_out & par_done_reg1054_out & par_done_reg1055_out & par_done_reg1056_out & par_done_reg1057_out & par_done_reg1058_out & par_done_reg1059_out & par_done_reg1060_out & par_done_reg1061_out & par_done_reg1062_out & par_done_reg1063_out & par_done_reg1064_out & par_done_reg1065_out & par_done_reg1066_out & par_done_reg1067_out & par_done_reg1068_out & par_done_reg1069_out & par_done_reg1070_out & par_done_reg1071_out & par_done_reg1072_out & par_done_reg1073_out & par_done_reg1074_out & par_done_reg1075_out & par_done_reg1076_out & par_done_reg1077_out & par_done_reg1078_out & par_done_reg1079_out & par_done_reg1080_out & par_done_reg1081_out & par_done_reg1082_out & par_done_reg1083_out & par_done_reg1084_out & par_done_reg1085_out & par_done_reg1086_out & par_done_reg1087_out & par_done_reg1088_out & par_done_reg1089_out & par_done_reg1090_out & par_done_reg1091_out & par_done_reg1092_out & par_done_reg1093_out & par_done_reg1094_out & par_done_reg1095_out & par_done_reg1096_out & par_done_reg1097_out & par_done_reg1098_out & par_done_reg1099_out & par_done_reg1100_out & par_done_reg1101_out & par_done_reg1102_out & par_done_reg1103_out & par_done_reg1104_out & par_done_reg1105_out & par_done_reg1106_out & par_done_reg1107_out & par_done_reg1108_out & par_done_reg1109_out & par_done_reg1110_out & par_done_reg1111_out & par_done_reg1112_out & par_done_reg1113_out & par_done_reg1114_out & par_done_reg1115_out & par_done_reg1116_out & par_done_reg1117_out & par_done_reg1118_out & par_done_reg1119_out & par_done_reg1120_out & par_done_reg1121_out & par_done_reg1122_out & par_done_reg1123_out & par_done_reg1124_out & par_done_reg1125_out & par_done_reg1126_out & par_done_reg1127_out & par_done_reg1128_out & par_done_reg1129_out & par_done_reg1130_out & par_done_reg1131_out & par_done_reg1132_out & par_done_reg1133_out & par_done_reg1134_out & par_done_reg1135_out & par_done_reg1136_out & par_done_reg1137_out & par_done_reg1138_out & par_done_reg1139_out & par_done_reg1140_out & par_done_reg1141_out & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_reset26_write_en = (par_done_reg1050_out & par_done_reg1051_out & par_done_reg1052_out & par_done_reg1053_out & par_done_reg1054_out & par_done_reg1055_out & par_done_reg1056_out & par_done_reg1057_out & par_done_reg1058_out & par_done_reg1059_out & par_done_reg1060_out & par_done_reg1061_out & par_done_reg1062_out & par_done_reg1063_out & par_done_reg1064_out & par_done_reg1065_out & par_done_reg1066_out & par_done_reg1067_out & par_done_reg1068_out & par_done_reg1069_out & par_done_reg1070_out & par_done_reg1071_out & par_done_reg1072_out & par_done_reg1073_out & par_done_reg1074_out & par_done_reg1075_out & par_done_reg1076_out & par_done_reg1077_out & par_done_reg1078_out & par_done_reg1079_out & par_done_reg1080_out & par_done_reg1081_out & par_done_reg1082_out & par_done_reg1083_out & par_done_reg1084_out & par_done_reg1085_out & par_done_reg1086_out & par_done_reg1087_out & par_done_reg1088_out & par_done_reg1089_out & par_done_reg1090_out & par_done_reg1091_out & par_done_reg1092_out & par_done_reg1093_out & par_done_reg1094_out & par_done_reg1095_out & par_done_reg1096_out & par_done_reg1097_out & par_done_reg1098_out & par_done_reg1099_out & par_done_reg1100_out & par_done_reg1101_out & par_done_reg1102_out & par_done_reg1103_out & par_done_reg1104_out & par_done_reg1105_out & par_done_reg1106_out & par_done_reg1107_out & par_done_reg1108_out & par_done_reg1109_out & par_done_reg1110_out & par_done_reg1111_out & par_done_reg1112_out & par_done_reg1113_out & par_done_reg1114_out & par_done_reg1115_out & par_done_reg1116_out & par_done_reg1117_out & par_done_reg1118_out & par_done_reg1119_out & par_done_reg1120_out & par_done_reg1121_out & par_done_reg1122_out & par_done_reg1123_out & par_done_reg1124_out & par_done_reg1125_out & par_done_reg1126_out & par_done_reg1127_out & par_done_reg1128_out & par_done_reg1129_out & par_done_reg1130_out & par_done_reg1131_out & par_done_reg1132_out & par_done_reg1133_out & par_done_reg1134_out & par_done_reg1135_out & par_done_reg1136_out & par_done_reg1137_out & par_done_reg1138_out & par_done_reg1139_out & par_done_reg1140_out & par_done_reg1141_out & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1050_in = par_reset26_out ? 1'd0 : (top_05_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1050_write_en = (top_05_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1051_in = par_reset26_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1051_write_en = (top_06_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1052_in = par_reset26_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1052_write_en = (top_07_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1053_in = par_reset26_out ? 1'd0 : (top_14_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1053_write_en = (top_14_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1054_in = par_reset26_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1054_write_en = (top_15_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1055_in = par_reset26_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1055_write_en = (top_16_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1056_in = par_reset26_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1056_write_en = (top_17_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1057_in = par_reset26_out ? 1'd0 : (top_23_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1057_write_en = (top_23_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1058_in = par_reset26_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1058_write_en = (top_24_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1059_in = par_reset26_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1059_write_en = (top_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1060_in = par_reset26_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1060_write_en = (top_26_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1061_in = par_reset26_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1061_write_en = (top_27_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1062_in = par_reset26_out ? 1'd0 : (top_32_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1062_write_en = (top_32_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1063_in = par_reset26_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1063_write_en = (top_33_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1064_in = par_reset26_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1064_write_en = (top_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1065_in = par_reset26_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1065_write_en = (top_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1066_in = par_reset26_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1066_write_en = (top_36_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1067_in = par_reset26_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1067_write_en = (top_37_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1068_in = par_reset26_out ? 1'd0 : (top_41_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1068_write_en = (top_41_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1069_in = par_reset26_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1069_write_en = (top_42_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1070_in = par_reset26_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1070_write_en = (top_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1071_in = par_reset26_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1071_write_en = (top_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1072_in = par_reset26_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1072_write_en = (top_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1073_in = par_reset26_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1073_write_en = (top_46_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1074_in = par_reset26_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1074_write_en = (top_47_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1075_in = par_reset26_out ? 1'd0 : (top_50_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1075_write_en = (top_50_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1076_in = par_reset26_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1076_write_en = (top_51_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1077_in = par_reset26_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1077_write_en = (top_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1078_in = par_reset26_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1078_write_en = (top_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1079_in = par_reset26_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1079_write_en = (top_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1080_in = par_reset26_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1080_write_en = (top_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1081_in = par_reset26_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1081_write_en = (top_56_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1082_in = par_reset26_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1082_write_en = (top_57_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1083_in = par_reset26_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1083_write_en = (top_60_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1084_in = par_reset26_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1084_write_en = (top_61_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1085_in = par_reset26_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1085_write_en = (top_62_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1086_in = par_reset26_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1086_write_en = (top_63_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1087_in = par_reset26_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1087_write_en = (top_64_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1088_in = par_reset26_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1088_write_en = (top_65_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1089_in = par_reset26_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1089_write_en = (top_66_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1090_in = par_reset26_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1090_write_en = (top_70_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1091_in = par_reset26_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1091_write_en = (top_71_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1092_in = par_reset26_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1092_write_en = (top_72_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1093_in = par_reset26_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1093_write_en = (top_73_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1094_in = par_reset26_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1094_write_en = (top_74_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1095_in = par_reset26_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1095_write_en = (top_75_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1096_in = par_reset26_out ? 1'd0 : (left_05_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1096_write_en = (left_05_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1097_in = par_reset26_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1097_write_en = (left_06_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1098_in = par_reset26_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1098_write_en = (left_07_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1099_in = par_reset26_out ? 1'd0 : (left_14_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1099_write_en = (left_14_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1100_in = par_reset26_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1100_write_en = (left_15_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1101_in = par_reset26_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1101_write_en = (left_16_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1102_in = par_reset26_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1102_write_en = (left_17_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1103_in = par_reset26_out ? 1'd0 : (left_23_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1103_write_en = (left_23_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1104_in = par_reset26_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1104_write_en = (left_24_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1105_in = par_reset26_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1105_write_en = (left_25_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1106_in = par_reset26_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1106_write_en = (left_26_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1107_in = par_reset26_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1107_write_en = (left_27_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1108_in = par_reset26_out ? 1'd0 : (left_32_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1108_write_en = (left_32_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1109_in = par_reset26_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1109_write_en = (left_33_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1110_in = par_reset26_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1110_write_en = (left_34_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1111_in = par_reset26_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1111_write_en = (left_35_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1112_in = par_reset26_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1112_write_en = (left_36_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1113_in = par_reset26_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1113_write_en = (left_37_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1114_in = par_reset26_out ? 1'd0 : (left_41_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1114_write_en = (left_41_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1115_in = par_reset26_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1115_write_en = (left_42_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1116_in = par_reset26_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1116_write_en = (left_43_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1117_in = par_reset26_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1117_write_en = (left_44_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1118_in = par_reset26_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1118_write_en = (left_45_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1119_in = par_reset26_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1119_write_en = (left_46_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1120_in = par_reset26_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1120_write_en = (left_47_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1121_in = par_reset26_out ? 1'd0 : (left_50_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1121_write_en = (left_50_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1122_in = par_reset26_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1122_write_en = (left_51_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1123_in = par_reset26_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1123_write_en = (left_52_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1124_in = par_reset26_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1124_write_en = (left_53_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1125_in = par_reset26_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1125_write_en = (left_54_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1126_in = par_reset26_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1126_write_en = (left_55_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1127_in = par_reset26_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1127_write_en = (left_56_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1128_in = par_reset26_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1128_write_en = (left_57_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1129_in = par_reset26_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1129_write_en = (left_60_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1130_in = par_reset26_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1130_write_en = (left_61_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1131_in = par_reset26_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1131_write_en = (left_62_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1132_in = par_reset26_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1132_write_en = (left_63_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1133_in = par_reset26_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1133_write_en = (left_64_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1134_in = par_reset26_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1134_write_en = (left_65_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1135_in = par_reset26_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1135_write_en = (left_66_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1136_in = par_reset26_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1136_write_en = (left_70_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1137_in = par_reset26_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1137_write_en = (left_71_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1138_in = par_reset26_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1138_write_en = (left_72_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1139_in = par_reset26_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1139_write_en = (left_73_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1140_in = par_reset26_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1140_write_en = (left_74_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_done_reg1141_in = par_reset26_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd26 & !par_reset26_out & go) ? 1'd1 : '0;
  assign par_done_reg1141_write_en = (left_75_read_done & fsm0_out == 32'd26 & !par_reset26_out & go | par_reset26_out) ? 1'd1 : '0;
  assign par_reset27_in = par_reset27_out ? 1'd0 : (par_done_reg1142_out & par_done_reg1143_out & par_done_reg1144_out & par_done_reg1145_out & par_done_reg1146_out & par_done_reg1147_out & par_done_reg1148_out & par_done_reg1149_out & par_done_reg1150_out & par_done_reg1151_out & par_done_reg1152_out & par_done_reg1153_out & par_done_reg1154_out & par_done_reg1155_out & par_done_reg1156_out & par_done_reg1157_out & par_done_reg1158_out & par_done_reg1159_out & par_done_reg1160_out & par_done_reg1161_out & par_done_reg1162_out & par_done_reg1163_out & par_done_reg1164_out & par_done_reg1165_out & par_done_reg1166_out & par_done_reg1167_out & par_done_reg1168_out & par_done_reg1169_out & par_done_reg1170_out & par_done_reg1171_out & par_done_reg1172_out & par_done_reg1173_out & par_done_reg1174_out & par_done_reg1175_out & par_done_reg1176_out & par_done_reg1177_out & par_done_reg1178_out & par_done_reg1179_out & par_done_reg1180_out & par_done_reg1181_out & par_done_reg1182_out & par_done_reg1183_out & par_done_reg1184_out & par_done_reg1185_out & par_done_reg1186_out & par_done_reg1187_out & par_done_reg1188_out & par_done_reg1189_out & par_done_reg1190_out & par_done_reg1191_out & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_reset27_write_en = (par_done_reg1142_out & par_done_reg1143_out & par_done_reg1144_out & par_done_reg1145_out & par_done_reg1146_out & par_done_reg1147_out & par_done_reg1148_out & par_done_reg1149_out & par_done_reg1150_out & par_done_reg1151_out & par_done_reg1152_out & par_done_reg1153_out & par_done_reg1154_out & par_done_reg1155_out & par_done_reg1156_out & par_done_reg1157_out & par_done_reg1158_out & par_done_reg1159_out & par_done_reg1160_out & par_done_reg1161_out & par_done_reg1162_out & par_done_reg1163_out & par_done_reg1164_out & par_done_reg1165_out & par_done_reg1166_out & par_done_reg1167_out & par_done_reg1168_out & par_done_reg1169_out & par_done_reg1170_out & par_done_reg1171_out & par_done_reg1172_out & par_done_reg1173_out & par_done_reg1174_out & par_done_reg1175_out & par_done_reg1176_out & par_done_reg1177_out & par_done_reg1178_out & par_done_reg1179_out & par_done_reg1180_out & par_done_reg1181_out & par_done_reg1182_out & par_done_reg1183_out & par_done_reg1184_out & par_done_reg1185_out & par_done_reg1186_out & par_done_reg1187_out & par_done_reg1188_out & par_done_reg1189_out & par_done_reg1190_out & par_done_reg1191_out & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1142_in = par_reset27_out ? 1'd0 : (t6_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1142_write_en = (t6_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1143_in = par_reset27_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1143_write_en = (t7_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1144_in = par_reset27_out ? 1'd0 : (l6_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1144_write_en = (l6_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1145_in = par_reset27_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1145_write_en = (l7_idx_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1146_in = par_reset27_out ? 1'd0 : (right_05_write_done & down_05_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1146_write_en = (right_05_write_done & down_05_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1147_in = par_reset27_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1147_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1148_in = par_reset27_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1148_write_en = (down_07_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1149_in = par_reset27_out ? 1'd0 : (right_14_write_done & down_14_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1149_write_en = (right_14_write_done & down_14_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1150_in = par_reset27_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1150_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1151_in = par_reset27_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1151_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1152_in = par_reset27_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1152_write_en = (down_17_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1153_in = par_reset27_out ? 1'd0 : (right_23_write_done & down_23_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1153_write_en = (right_23_write_done & down_23_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1154_in = par_reset27_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1154_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1155_in = par_reset27_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1155_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1156_in = par_reset27_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1156_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1157_in = par_reset27_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1157_write_en = (down_27_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1158_in = par_reset27_out ? 1'd0 : (right_32_write_done & down_32_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1158_write_en = (right_32_write_done & down_32_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1159_in = par_reset27_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1159_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1160_in = par_reset27_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1160_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1161_in = par_reset27_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1161_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1162_in = par_reset27_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1162_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1163_in = par_reset27_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1163_write_en = (down_37_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1164_in = par_reset27_out ? 1'd0 : (right_41_write_done & down_41_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1164_write_en = (right_41_write_done & down_41_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1165_in = par_reset27_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1165_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1166_in = par_reset27_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1166_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1167_in = par_reset27_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1167_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1168_in = par_reset27_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1168_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1169_in = par_reset27_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1169_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1170_in = par_reset27_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1170_write_en = (down_47_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1171_in = par_reset27_out ? 1'd0 : (right_50_write_done & down_50_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1171_write_en = (right_50_write_done & down_50_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1172_in = par_reset27_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1172_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1173_in = par_reset27_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1173_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1174_in = par_reset27_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1174_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1175_in = par_reset27_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1175_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1176_in = par_reset27_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1176_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1177_in = par_reset27_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1177_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1178_in = par_reset27_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1178_write_en = (down_57_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1179_in = par_reset27_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1179_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1180_in = par_reset27_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1180_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1181_in = par_reset27_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1181_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1182_in = par_reset27_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1182_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1183_in = par_reset27_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1183_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1184_in = par_reset27_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1184_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1185_in = par_reset27_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1185_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1186_in = par_reset27_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1186_write_en = (right_70_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1187_in = par_reset27_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1187_write_en = (right_71_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1188_in = par_reset27_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1188_write_en = (right_72_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1189_in = par_reset27_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1189_write_en = (right_73_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1190_in = par_reset27_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1190_write_en = (right_74_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_done_reg1191_in = par_reset27_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd27 & !par_reset27_out & go) ? 1'd1 : '0;
  assign par_done_reg1191_write_en = (right_75_write_done & fsm0_out == 32'd27 & !par_reset27_out & go | par_reset27_out) ? 1'd1 : '0;
  assign par_reset28_in = par_reset28_out ? 1'd0 : (par_done_reg1192_out & par_done_reg1193_out & par_done_reg1194_out & par_done_reg1195_out & par_done_reg1196_out & par_done_reg1197_out & par_done_reg1198_out & par_done_reg1199_out & par_done_reg1200_out & par_done_reg1201_out & par_done_reg1202_out & par_done_reg1203_out & par_done_reg1204_out & par_done_reg1205_out & par_done_reg1206_out & par_done_reg1207_out & par_done_reg1208_out & par_done_reg1209_out & par_done_reg1210_out & par_done_reg1211_out & par_done_reg1212_out & par_done_reg1213_out & par_done_reg1214_out & par_done_reg1215_out & par_done_reg1216_out & par_done_reg1217_out & par_done_reg1218_out & par_done_reg1219_out & par_done_reg1220_out & par_done_reg1221_out & par_done_reg1222_out & par_done_reg1223_out & par_done_reg1224_out & par_done_reg1225_out & par_done_reg1226_out & par_done_reg1227_out & par_done_reg1228_out & par_done_reg1229_out & par_done_reg1230_out & par_done_reg1231_out & par_done_reg1232_out & par_done_reg1233_out & par_done_reg1234_out & par_done_reg1235_out & par_done_reg1236_out & par_done_reg1237_out & par_done_reg1238_out & par_done_reg1239_out & par_done_reg1240_out & par_done_reg1241_out & par_done_reg1242_out & par_done_reg1243_out & par_done_reg1244_out & par_done_reg1245_out & par_done_reg1246_out & par_done_reg1247_out & par_done_reg1248_out & par_done_reg1249_out & par_done_reg1250_out & par_done_reg1251_out & par_done_reg1252_out & par_done_reg1253_out & par_done_reg1254_out & par_done_reg1255_out & par_done_reg1256_out & par_done_reg1257_out & par_done_reg1258_out & par_done_reg1259_out & par_done_reg1260_out & par_done_reg1261_out & par_done_reg1262_out & par_done_reg1263_out & par_done_reg1264_out & par_done_reg1265_out & par_done_reg1266_out & par_done_reg1267_out & par_done_reg1268_out & par_done_reg1269_out & par_done_reg1270_out & par_done_reg1271_out & par_done_reg1272_out & par_done_reg1273_out & par_done_reg1274_out & par_done_reg1275_out & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_reset28_write_en = (par_done_reg1192_out & par_done_reg1193_out & par_done_reg1194_out & par_done_reg1195_out & par_done_reg1196_out & par_done_reg1197_out & par_done_reg1198_out & par_done_reg1199_out & par_done_reg1200_out & par_done_reg1201_out & par_done_reg1202_out & par_done_reg1203_out & par_done_reg1204_out & par_done_reg1205_out & par_done_reg1206_out & par_done_reg1207_out & par_done_reg1208_out & par_done_reg1209_out & par_done_reg1210_out & par_done_reg1211_out & par_done_reg1212_out & par_done_reg1213_out & par_done_reg1214_out & par_done_reg1215_out & par_done_reg1216_out & par_done_reg1217_out & par_done_reg1218_out & par_done_reg1219_out & par_done_reg1220_out & par_done_reg1221_out & par_done_reg1222_out & par_done_reg1223_out & par_done_reg1224_out & par_done_reg1225_out & par_done_reg1226_out & par_done_reg1227_out & par_done_reg1228_out & par_done_reg1229_out & par_done_reg1230_out & par_done_reg1231_out & par_done_reg1232_out & par_done_reg1233_out & par_done_reg1234_out & par_done_reg1235_out & par_done_reg1236_out & par_done_reg1237_out & par_done_reg1238_out & par_done_reg1239_out & par_done_reg1240_out & par_done_reg1241_out & par_done_reg1242_out & par_done_reg1243_out & par_done_reg1244_out & par_done_reg1245_out & par_done_reg1246_out & par_done_reg1247_out & par_done_reg1248_out & par_done_reg1249_out & par_done_reg1250_out & par_done_reg1251_out & par_done_reg1252_out & par_done_reg1253_out & par_done_reg1254_out & par_done_reg1255_out & par_done_reg1256_out & par_done_reg1257_out & par_done_reg1258_out & par_done_reg1259_out & par_done_reg1260_out & par_done_reg1261_out & par_done_reg1262_out & par_done_reg1263_out & par_done_reg1264_out & par_done_reg1265_out & par_done_reg1266_out & par_done_reg1267_out & par_done_reg1268_out & par_done_reg1269_out & par_done_reg1270_out & par_done_reg1271_out & par_done_reg1272_out & par_done_reg1273_out & par_done_reg1274_out & par_done_reg1275_out & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1192_in = par_reset28_out ? 1'd0 : (top_06_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1192_write_en = (top_06_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1193_in = par_reset28_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1193_write_en = (top_07_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1194_in = par_reset28_out ? 1'd0 : (top_15_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1194_write_en = (top_15_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1195_in = par_reset28_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1195_write_en = (top_16_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1196_in = par_reset28_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1196_write_en = (top_17_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1197_in = par_reset28_out ? 1'd0 : (top_24_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1197_write_en = (top_24_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1198_in = par_reset28_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1198_write_en = (top_25_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1199_in = par_reset28_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1199_write_en = (top_26_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1200_in = par_reset28_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1200_write_en = (top_27_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1201_in = par_reset28_out ? 1'd0 : (top_33_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1201_write_en = (top_33_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1202_in = par_reset28_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1202_write_en = (top_34_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1203_in = par_reset28_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1203_write_en = (top_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1204_in = par_reset28_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1204_write_en = (top_36_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1205_in = par_reset28_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1205_write_en = (top_37_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1206_in = par_reset28_out ? 1'd0 : (top_42_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1206_write_en = (top_42_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1207_in = par_reset28_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1207_write_en = (top_43_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1208_in = par_reset28_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1208_write_en = (top_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1209_in = par_reset28_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1209_write_en = (top_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1210_in = par_reset28_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1210_write_en = (top_46_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1211_in = par_reset28_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1211_write_en = (top_47_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1212_in = par_reset28_out ? 1'd0 : (top_51_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1212_write_en = (top_51_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1213_in = par_reset28_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1213_write_en = (top_52_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1214_in = par_reset28_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1214_write_en = (top_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1215_in = par_reset28_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1215_write_en = (top_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1216_in = par_reset28_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1216_write_en = (top_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1217_in = par_reset28_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1217_write_en = (top_56_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1218_in = par_reset28_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1218_write_en = (top_57_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1219_in = par_reset28_out ? 1'd0 : (top_60_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1219_write_en = (top_60_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1220_in = par_reset28_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1220_write_en = (top_61_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1221_in = par_reset28_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1221_write_en = (top_62_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1222_in = par_reset28_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1222_write_en = (top_63_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1223_in = par_reset28_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1223_write_en = (top_64_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1224_in = par_reset28_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1224_write_en = (top_65_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1225_in = par_reset28_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1225_write_en = (top_66_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1226_in = par_reset28_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1226_write_en = (top_67_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1227_in = par_reset28_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1227_write_en = (top_70_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1228_in = par_reset28_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1228_write_en = (top_71_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1229_in = par_reset28_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1229_write_en = (top_72_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1230_in = par_reset28_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1230_write_en = (top_73_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1231_in = par_reset28_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1231_write_en = (top_74_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1232_in = par_reset28_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1232_write_en = (top_75_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1233_in = par_reset28_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1233_write_en = (top_76_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1234_in = par_reset28_out ? 1'd0 : (left_06_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1234_write_en = (left_06_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1235_in = par_reset28_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1235_write_en = (left_07_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1236_in = par_reset28_out ? 1'd0 : (left_15_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1236_write_en = (left_15_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1237_in = par_reset28_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1237_write_en = (left_16_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1238_in = par_reset28_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1238_write_en = (left_17_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1239_in = par_reset28_out ? 1'd0 : (left_24_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1239_write_en = (left_24_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1240_in = par_reset28_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1240_write_en = (left_25_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1241_in = par_reset28_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1241_write_en = (left_26_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1242_in = par_reset28_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1242_write_en = (left_27_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1243_in = par_reset28_out ? 1'd0 : (left_33_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1243_write_en = (left_33_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1244_in = par_reset28_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1244_write_en = (left_34_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1245_in = par_reset28_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1245_write_en = (left_35_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1246_in = par_reset28_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1246_write_en = (left_36_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1247_in = par_reset28_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1247_write_en = (left_37_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1248_in = par_reset28_out ? 1'd0 : (left_42_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1248_write_en = (left_42_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1249_in = par_reset28_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1249_write_en = (left_43_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1250_in = par_reset28_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1250_write_en = (left_44_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1251_in = par_reset28_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1251_write_en = (left_45_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1252_in = par_reset28_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1252_write_en = (left_46_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1253_in = par_reset28_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1253_write_en = (left_47_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1254_in = par_reset28_out ? 1'd0 : (left_51_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1254_write_en = (left_51_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1255_in = par_reset28_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1255_write_en = (left_52_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1256_in = par_reset28_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1256_write_en = (left_53_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1257_in = par_reset28_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1257_write_en = (left_54_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1258_in = par_reset28_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1258_write_en = (left_55_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1259_in = par_reset28_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1259_write_en = (left_56_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1260_in = par_reset28_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1260_write_en = (left_57_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1261_in = par_reset28_out ? 1'd0 : (left_60_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1261_write_en = (left_60_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1262_in = par_reset28_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1262_write_en = (left_61_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1263_in = par_reset28_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1263_write_en = (left_62_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1264_in = par_reset28_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1264_write_en = (left_63_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1265_in = par_reset28_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1265_write_en = (left_64_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1266_in = par_reset28_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1266_write_en = (left_65_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1267_in = par_reset28_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1267_write_en = (left_66_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1268_in = par_reset28_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1268_write_en = (left_67_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1269_in = par_reset28_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1269_write_en = (left_70_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1270_in = par_reset28_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1270_write_en = (left_71_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1271_in = par_reset28_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1271_write_en = (left_72_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1272_in = par_reset28_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1272_write_en = (left_73_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1273_in = par_reset28_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1273_write_en = (left_74_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1274_in = par_reset28_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1274_write_en = (left_75_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_done_reg1275_in = par_reset28_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd28 & !par_reset28_out & go) ? 1'd1 : '0;
  assign par_done_reg1275_write_en = (left_76_read_done & fsm0_out == 32'd28 & !par_reset28_out & go | par_reset28_out) ? 1'd1 : '0;
  assign par_reset29_in = par_reset29_out ? 1'd0 : (par_done_reg1276_out & par_done_reg1277_out & par_done_reg1278_out & par_done_reg1279_out & par_done_reg1280_out & par_done_reg1281_out & par_done_reg1282_out & par_done_reg1283_out & par_done_reg1284_out & par_done_reg1285_out & par_done_reg1286_out & par_done_reg1287_out & par_done_reg1288_out & par_done_reg1289_out & par_done_reg1290_out & par_done_reg1291_out & par_done_reg1292_out & par_done_reg1293_out & par_done_reg1294_out & par_done_reg1295_out & par_done_reg1296_out & par_done_reg1297_out & par_done_reg1298_out & par_done_reg1299_out & par_done_reg1300_out & par_done_reg1301_out & par_done_reg1302_out & par_done_reg1303_out & par_done_reg1304_out & par_done_reg1305_out & par_done_reg1306_out & par_done_reg1307_out & par_done_reg1308_out & par_done_reg1309_out & par_done_reg1310_out & par_done_reg1311_out & par_done_reg1312_out & par_done_reg1313_out & par_done_reg1314_out & par_done_reg1315_out & par_done_reg1316_out & par_done_reg1317_out & par_done_reg1318_out & par_done_reg1319_out & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_reset29_write_en = (par_done_reg1276_out & par_done_reg1277_out & par_done_reg1278_out & par_done_reg1279_out & par_done_reg1280_out & par_done_reg1281_out & par_done_reg1282_out & par_done_reg1283_out & par_done_reg1284_out & par_done_reg1285_out & par_done_reg1286_out & par_done_reg1287_out & par_done_reg1288_out & par_done_reg1289_out & par_done_reg1290_out & par_done_reg1291_out & par_done_reg1292_out & par_done_reg1293_out & par_done_reg1294_out & par_done_reg1295_out & par_done_reg1296_out & par_done_reg1297_out & par_done_reg1298_out & par_done_reg1299_out & par_done_reg1300_out & par_done_reg1301_out & par_done_reg1302_out & par_done_reg1303_out & par_done_reg1304_out & par_done_reg1305_out & par_done_reg1306_out & par_done_reg1307_out & par_done_reg1308_out & par_done_reg1309_out & par_done_reg1310_out & par_done_reg1311_out & par_done_reg1312_out & par_done_reg1313_out & par_done_reg1314_out & par_done_reg1315_out & par_done_reg1316_out & par_done_reg1317_out & par_done_reg1318_out & par_done_reg1319_out & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1276_in = par_reset29_out ? 1'd0 : (t7_idx_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1276_write_en = (t7_idx_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1277_in = par_reset29_out ? 1'd0 : (l7_idx_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1277_write_en = (l7_idx_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1278_in = par_reset29_out ? 1'd0 : (right_06_write_done & down_06_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1278_write_en = (right_06_write_done & down_06_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1279_in = par_reset29_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1279_write_en = (down_07_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1280_in = par_reset29_out ? 1'd0 : (right_15_write_done & down_15_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1280_write_en = (right_15_write_done & down_15_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1281_in = par_reset29_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1281_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1282_in = par_reset29_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1282_write_en = (down_17_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1283_in = par_reset29_out ? 1'd0 : (right_24_write_done & down_24_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1283_write_en = (right_24_write_done & down_24_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1284_in = par_reset29_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1284_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1285_in = par_reset29_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1285_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1286_in = par_reset29_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1286_write_en = (down_27_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1287_in = par_reset29_out ? 1'd0 : (right_33_write_done & down_33_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1287_write_en = (right_33_write_done & down_33_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1288_in = par_reset29_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1288_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1289_in = par_reset29_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1289_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1290_in = par_reset29_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1290_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1291_in = par_reset29_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1291_write_en = (down_37_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1292_in = par_reset29_out ? 1'd0 : (right_42_write_done & down_42_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1292_write_en = (right_42_write_done & down_42_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1293_in = par_reset29_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1293_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1294_in = par_reset29_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1294_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1295_in = par_reset29_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1295_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1296_in = par_reset29_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1296_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1297_in = par_reset29_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1297_write_en = (down_47_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1298_in = par_reset29_out ? 1'd0 : (right_51_write_done & down_51_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1298_write_en = (right_51_write_done & down_51_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1299_in = par_reset29_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1299_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1300_in = par_reset29_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1300_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1301_in = par_reset29_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1301_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1302_in = par_reset29_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1302_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1303_in = par_reset29_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1303_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1304_in = par_reset29_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1304_write_en = (down_57_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1305_in = par_reset29_out ? 1'd0 : (right_60_write_done & down_60_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1305_write_en = (right_60_write_done & down_60_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1306_in = par_reset29_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1306_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1307_in = par_reset29_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1307_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1308_in = par_reset29_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1308_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1309_in = par_reset29_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1309_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1310_in = par_reset29_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1310_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1311_in = par_reset29_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1311_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1312_in = par_reset29_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1312_write_en = (down_67_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1313_in = par_reset29_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1313_write_en = (right_70_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1314_in = par_reset29_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1314_write_en = (right_71_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1315_in = par_reset29_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1315_write_en = (right_72_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1316_in = par_reset29_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1316_write_en = (right_73_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1317_in = par_reset29_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1317_write_en = (right_74_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1318_in = par_reset29_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1318_write_en = (right_75_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_done_reg1319_in = par_reset29_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd29 & !par_reset29_out & go) ? 1'd1 : '0;
  assign par_done_reg1319_write_en = (right_76_write_done & fsm0_out == 32'd29 & !par_reset29_out & go | par_reset29_out) ? 1'd1 : '0;
  assign par_reset30_in = par_reset30_out ? 1'd0 : (par_done_reg1320_out & par_done_reg1321_out & par_done_reg1322_out & par_done_reg1323_out & par_done_reg1324_out & par_done_reg1325_out & par_done_reg1326_out & par_done_reg1327_out & par_done_reg1328_out & par_done_reg1329_out & par_done_reg1330_out & par_done_reg1331_out & par_done_reg1332_out & par_done_reg1333_out & par_done_reg1334_out & par_done_reg1335_out & par_done_reg1336_out & par_done_reg1337_out & par_done_reg1338_out & par_done_reg1339_out & par_done_reg1340_out & par_done_reg1341_out & par_done_reg1342_out & par_done_reg1343_out & par_done_reg1344_out & par_done_reg1345_out & par_done_reg1346_out & par_done_reg1347_out & par_done_reg1348_out & par_done_reg1349_out & par_done_reg1350_out & par_done_reg1351_out & par_done_reg1352_out & par_done_reg1353_out & par_done_reg1354_out & par_done_reg1355_out & par_done_reg1356_out & par_done_reg1357_out & par_done_reg1358_out & par_done_reg1359_out & par_done_reg1360_out & par_done_reg1361_out & par_done_reg1362_out & par_done_reg1363_out & par_done_reg1364_out & par_done_reg1365_out & par_done_reg1366_out & par_done_reg1367_out & par_done_reg1368_out & par_done_reg1369_out & par_done_reg1370_out & par_done_reg1371_out & par_done_reg1372_out & par_done_reg1373_out & par_done_reg1374_out & par_done_reg1375_out & par_done_reg1376_out & par_done_reg1377_out & par_done_reg1378_out & par_done_reg1379_out & par_done_reg1380_out & par_done_reg1381_out & par_done_reg1382_out & par_done_reg1383_out & par_done_reg1384_out & par_done_reg1385_out & par_done_reg1386_out & par_done_reg1387_out & par_done_reg1388_out & par_done_reg1389_out & par_done_reg1390_out & par_done_reg1391_out & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_reset30_write_en = (par_done_reg1320_out & par_done_reg1321_out & par_done_reg1322_out & par_done_reg1323_out & par_done_reg1324_out & par_done_reg1325_out & par_done_reg1326_out & par_done_reg1327_out & par_done_reg1328_out & par_done_reg1329_out & par_done_reg1330_out & par_done_reg1331_out & par_done_reg1332_out & par_done_reg1333_out & par_done_reg1334_out & par_done_reg1335_out & par_done_reg1336_out & par_done_reg1337_out & par_done_reg1338_out & par_done_reg1339_out & par_done_reg1340_out & par_done_reg1341_out & par_done_reg1342_out & par_done_reg1343_out & par_done_reg1344_out & par_done_reg1345_out & par_done_reg1346_out & par_done_reg1347_out & par_done_reg1348_out & par_done_reg1349_out & par_done_reg1350_out & par_done_reg1351_out & par_done_reg1352_out & par_done_reg1353_out & par_done_reg1354_out & par_done_reg1355_out & par_done_reg1356_out & par_done_reg1357_out & par_done_reg1358_out & par_done_reg1359_out & par_done_reg1360_out & par_done_reg1361_out & par_done_reg1362_out & par_done_reg1363_out & par_done_reg1364_out & par_done_reg1365_out & par_done_reg1366_out & par_done_reg1367_out & par_done_reg1368_out & par_done_reg1369_out & par_done_reg1370_out & par_done_reg1371_out & par_done_reg1372_out & par_done_reg1373_out & par_done_reg1374_out & par_done_reg1375_out & par_done_reg1376_out & par_done_reg1377_out & par_done_reg1378_out & par_done_reg1379_out & par_done_reg1380_out & par_done_reg1381_out & par_done_reg1382_out & par_done_reg1383_out & par_done_reg1384_out & par_done_reg1385_out & par_done_reg1386_out & par_done_reg1387_out & par_done_reg1388_out & par_done_reg1389_out & par_done_reg1390_out & par_done_reg1391_out & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1320_in = par_reset30_out ? 1'd0 : (top_07_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1320_write_en = (top_07_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1321_in = par_reset30_out ? 1'd0 : (top_16_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1321_write_en = (top_16_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1322_in = par_reset30_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1322_write_en = (top_17_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1323_in = par_reset30_out ? 1'd0 : (top_25_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1323_write_en = (top_25_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1324_in = par_reset30_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1324_write_en = (top_26_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1325_in = par_reset30_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1325_write_en = (top_27_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1326_in = par_reset30_out ? 1'd0 : (top_34_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1326_write_en = (top_34_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1327_in = par_reset30_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1327_write_en = (top_35_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1328_in = par_reset30_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1328_write_en = (top_36_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1329_in = par_reset30_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1329_write_en = (top_37_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1330_in = par_reset30_out ? 1'd0 : (top_43_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1330_write_en = (top_43_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1331_in = par_reset30_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1331_write_en = (top_44_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1332_in = par_reset30_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1332_write_en = (top_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1333_in = par_reset30_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1333_write_en = (top_46_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1334_in = par_reset30_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1334_write_en = (top_47_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1335_in = par_reset30_out ? 1'd0 : (top_52_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1335_write_en = (top_52_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1336_in = par_reset30_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1336_write_en = (top_53_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1337_in = par_reset30_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1337_write_en = (top_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1338_in = par_reset30_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1338_write_en = (top_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1339_in = par_reset30_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1339_write_en = (top_56_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1340_in = par_reset30_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1340_write_en = (top_57_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1341_in = par_reset30_out ? 1'd0 : (top_61_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1341_write_en = (top_61_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1342_in = par_reset30_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1342_write_en = (top_62_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1343_in = par_reset30_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1343_write_en = (top_63_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1344_in = par_reset30_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1344_write_en = (top_64_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1345_in = par_reset30_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1345_write_en = (top_65_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1346_in = par_reset30_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1346_write_en = (top_66_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1347_in = par_reset30_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1347_write_en = (top_67_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1348_in = par_reset30_out ? 1'd0 : (top_70_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1348_write_en = (top_70_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1349_in = par_reset30_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1349_write_en = (top_71_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1350_in = par_reset30_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1350_write_en = (top_72_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1351_in = par_reset30_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1351_write_en = (top_73_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1352_in = par_reset30_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1352_write_en = (top_74_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1353_in = par_reset30_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1353_write_en = (top_75_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1354_in = par_reset30_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1354_write_en = (top_76_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1355_in = par_reset30_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1355_write_en = (top_77_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1356_in = par_reset30_out ? 1'd0 : (left_07_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1356_write_en = (left_07_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1357_in = par_reset30_out ? 1'd0 : (left_16_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1357_write_en = (left_16_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1358_in = par_reset30_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1358_write_en = (left_17_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1359_in = par_reset30_out ? 1'd0 : (left_25_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1359_write_en = (left_25_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1360_in = par_reset30_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1360_write_en = (left_26_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1361_in = par_reset30_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1361_write_en = (left_27_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1362_in = par_reset30_out ? 1'd0 : (left_34_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1362_write_en = (left_34_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1363_in = par_reset30_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1363_write_en = (left_35_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1364_in = par_reset30_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1364_write_en = (left_36_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1365_in = par_reset30_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1365_write_en = (left_37_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1366_in = par_reset30_out ? 1'd0 : (left_43_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1366_write_en = (left_43_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1367_in = par_reset30_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1367_write_en = (left_44_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1368_in = par_reset30_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1368_write_en = (left_45_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1369_in = par_reset30_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1369_write_en = (left_46_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1370_in = par_reset30_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1370_write_en = (left_47_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1371_in = par_reset30_out ? 1'd0 : (left_52_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1371_write_en = (left_52_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1372_in = par_reset30_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1372_write_en = (left_53_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1373_in = par_reset30_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1373_write_en = (left_54_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1374_in = par_reset30_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1374_write_en = (left_55_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1375_in = par_reset30_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1375_write_en = (left_56_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1376_in = par_reset30_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1376_write_en = (left_57_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1377_in = par_reset30_out ? 1'd0 : (left_61_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1377_write_en = (left_61_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1378_in = par_reset30_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1378_write_en = (left_62_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1379_in = par_reset30_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1379_write_en = (left_63_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1380_in = par_reset30_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1380_write_en = (left_64_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1381_in = par_reset30_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1381_write_en = (left_65_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1382_in = par_reset30_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1382_write_en = (left_66_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1383_in = par_reset30_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1383_write_en = (left_67_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1384_in = par_reset30_out ? 1'd0 : (left_70_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1384_write_en = (left_70_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1385_in = par_reset30_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1385_write_en = (left_71_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1386_in = par_reset30_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1386_write_en = (left_72_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1387_in = par_reset30_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1387_write_en = (left_73_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1388_in = par_reset30_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1388_write_en = (left_74_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1389_in = par_reset30_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1389_write_en = (left_75_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1390_in = par_reset30_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1390_write_en = (left_76_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_done_reg1391_in = par_reset30_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd30 & !par_reset30_out & go) ? 1'd1 : '0;
  assign par_done_reg1391_write_en = (left_77_read_done & fsm0_out == 32'd30 & !par_reset30_out & go | par_reset30_out) ? 1'd1 : '0;
  assign par_reset31_in = par_reset31_out ? 1'd0 : (par_done_reg1392_out & par_done_reg1393_out & par_done_reg1394_out & par_done_reg1395_out & par_done_reg1396_out & par_done_reg1397_out & par_done_reg1398_out & par_done_reg1399_out & par_done_reg1400_out & par_done_reg1401_out & par_done_reg1402_out & par_done_reg1403_out & par_done_reg1404_out & par_done_reg1405_out & par_done_reg1406_out & par_done_reg1407_out & par_done_reg1408_out & par_done_reg1409_out & par_done_reg1410_out & par_done_reg1411_out & par_done_reg1412_out & par_done_reg1413_out & par_done_reg1414_out & par_done_reg1415_out & par_done_reg1416_out & par_done_reg1417_out & par_done_reg1418_out & par_done_reg1419_out & par_done_reg1420_out & par_done_reg1421_out & par_done_reg1422_out & par_done_reg1423_out & par_done_reg1424_out & par_done_reg1425_out & par_done_reg1426_out & par_done_reg1427_out & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_reset31_write_en = (par_done_reg1392_out & par_done_reg1393_out & par_done_reg1394_out & par_done_reg1395_out & par_done_reg1396_out & par_done_reg1397_out & par_done_reg1398_out & par_done_reg1399_out & par_done_reg1400_out & par_done_reg1401_out & par_done_reg1402_out & par_done_reg1403_out & par_done_reg1404_out & par_done_reg1405_out & par_done_reg1406_out & par_done_reg1407_out & par_done_reg1408_out & par_done_reg1409_out & par_done_reg1410_out & par_done_reg1411_out & par_done_reg1412_out & par_done_reg1413_out & par_done_reg1414_out & par_done_reg1415_out & par_done_reg1416_out & par_done_reg1417_out & par_done_reg1418_out & par_done_reg1419_out & par_done_reg1420_out & par_done_reg1421_out & par_done_reg1422_out & par_done_reg1423_out & par_done_reg1424_out & par_done_reg1425_out & par_done_reg1426_out & par_done_reg1427_out & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1392_in = par_reset31_out ? 1'd0 : (down_07_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1392_write_en = (down_07_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1393_in = par_reset31_out ? 1'd0 : (right_16_write_done & down_16_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1393_write_en = (right_16_write_done & down_16_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1394_in = par_reset31_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1394_write_en = (down_17_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1395_in = par_reset31_out ? 1'd0 : (right_25_write_done & down_25_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1395_write_en = (right_25_write_done & down_25_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1396_in = par_reset31_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1396_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1397_in = par_reset31_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1397_write_en = (down_27_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1398_in = par_reset31_out ? 1'd0 : (right_34_write_done & down_34_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1398_write_en = (right_34_write_done & down_34_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1399_in = par_reset31_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1399_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1400_in = par_reset31_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1400_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1401_in = par_reset31_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1401_write_en = (down_37_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1402_in = par_reset31_out ? 1'd0 : (right_43_write_done & down_43_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1402_write_en = (right_43_write_done & down_43_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1403_in = par_reset31_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1403_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1404_in = par_reset31_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1404_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1405_in = par_reset31_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1405_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1406_in = par_reset31_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1406_write_en = (down_47_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1407_in = par_reset31_out ? 1'd0 : (right_52_write_done & down_52_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1407_write_en = (right_52_write_done & down_52_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1408_in = par_reset31_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1408_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1409_in = par_reset31_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1409_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1410_in = par_reset31_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1410_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1411_in = par_reset31_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1411_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1412_in = par_reset31_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1412_write_en = (down_57_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1413_in = par_reset31_out ? 1'd0 : (right_61_write_done & down_61_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1413_write_en = (right_61_write_done & down_61_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1414_in = par_reset31_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1414_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1415_in = par_reset31_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1415_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1416_in = par_reset31_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1416_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1417_in = par_reset31_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1417_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1418_in = par_reset31_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1418_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1419_in = par_reset31_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1419_write_en = (down_67_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1420_in = par_reset31_out ? 1'd0 : (right_70_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1420_write_en = (right_70_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1421_in = par_reset31_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1421_write_en = (right_71_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1422_in = par_reset31_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1422_write_en = (right_72_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1423_in = par_reset31_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1423_write_en = (right_73_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1424_in = par_reset31_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1424_write_en = (right_74_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1425_in = par_reset31_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1425_write_en = (right_75_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1426_in = par_reset31_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1426_write_en = (right_76_write_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_done_reg1427_in = par_reset31_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd31 & !par_reset31_out & go) ? 1'd1 : '0;
  assign par_done_reg1427_write_en = (pe_77_done & fsm0_out == 32'd31 & !par_reset31_out & go | par_reset31_out) ? 1'd1 : '0;
  assign par_reset32_in = par_reset32_out ? 1'd0 : (par_done_reg1428_out & par_done_reg1429_out & par_done_reg1430_out & par_done_reg1431_out & par_done_reg1432_out & par_done_reg1433_out & par_done_reg1434_out & par_done_reg1435_out & par_done_reg1436_out & par_done_reg1437_out & par_done_reg1438_out & par_done_reg1439_out & par_done_reg1440_out & par_done_reg1441_out & par_done_reg1442_out & par_done_reg1443_out & par_done_reg1444_out & par_done_reg1445_out & par_done_reg1446_out & par_done_reg1447_out & par_done_reg1448_out & par_done_reg1449_out & par_done_reg1450_out & par_done_reg1451_out & par_done_reg1452_out & par_done_reg1453_out & par_done_reg1454_out & par_done_reg1455_out & par_done_reg1456_out & par_done_reg1457_out & par_done_reg1458_out & par_done_reg1459_out & par_done_reg1460_out & par_done_reg1461_out & par_done_reg1462_out & par_done_reg1463_out & par_done_reg1464_out & par_done_reg1465_out & par_done_reg1466_out & par_done_reg1467_out & par_done_reg1468_out & par_done_reg1469_out & par_done_reg1470_out & par_done_reg1471_out & par_done_reg1472_out & par_done_reg1473_out & par_done_reg1474_out & par_done_reg1475_out & par_done_reg1476_out & par_done_reg1477_out & par_done_reg1478_out & par_done_reg1479_out & par_done_reg1480_out & par_done_reg1481_out & par_done_reg1482_out & par_done_reg1483_out & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_reset32_write_en = (par_done_reg1428_out & par_done_reg1429_out & par_done_reg1430_out & par_done_reg1431_out & par_done_reg1432_out & par_done_reg1433_out & par_done_reg1434_out & par_done_reg1435_out & par_done_reg1436_out & par_done_reg1437_out & par_done_reg1438_out & par_done_reg1439_out & par_done_reg1440_out & par_done_reg1441_out & par_done_reg1442_out & par_done_reg1443_out & par_done_reg1444_out & par_done_reg1445_out & par_done_reg1446_out & par_done_reg1447_out & par_done_reg1448_out & par_done_reg1449_out & par_done_reg1450_out & par_done_reg1451_out & par_done_reg1452_out & par_done_reg1453_out & par_done_reg1454_out & par_done_reg1455_out & par_done_reg1456_out & par_done_reg1457_out & par_done_reg1458_out & par_done_reg1459_out & par_done_reg1460_out & par_done_reg1461_out & par_done_reg1462_out & par_done_reg1463_out & par_done_reg1464_out & par_done_reg1465_out & par_done_reg1466_out & par_done_reg1467_out & par_done_reg1468_out & par_done_reg1469_out & par_done_reg1470_out & par_done_reg1471_out & par_done_reg1472_out & par_done_reg1473_out & par_done_reg1474_out & par_done_reg1475_out & par_done_reg1476_out & par_done_reg1477_out & par_done_reg1478_out & par_done_reg1479_out & par_done_reg1480_out & par_done_reg1481_out & par_done_reg1482_out & par_done_reg1483_out & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1428_in = par_reset32_out ? 1'd0 : (top_17_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1428_write_en = (top_17_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1429_in = par_reset32_out ? 1'd0 : (top_26_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1429_write_en = (top_26_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1430_in = par_reset32_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1430_write_en = (top_27_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1431_in = par_reset32_out ? 1'd0 : (top_35_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1431_write_en = (top_35_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1432_in = par_reset32_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1432_write_en = (top_36_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1433_in = par_reset32_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1433_write_en = (top_37_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1434_in = par_reset32_out ? 1'd0 : (top_44_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1434_write_en = (top_44_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1435_in = par_reset32_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1435_write_en = (top_45_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1436_in = par_reset32_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1436_write_en = (top_46_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1437_in = par_reset32_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1437_write_en = (top_47_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1438_in = par_reset32_out ? 1'd0 : (top_53_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1438_write_en = (top_53_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1439_in = par_reset32_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1439_write_en = (top_54_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1440_in = par_reset32_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1440_write_en = (top_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1441_in = par_reset32_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1441_write_en = (top_56_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1442_in = par_reset32_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1442_write_en = (top_57_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1443_in = par_reset32_out ? 1'd0 : (top_62_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1443_write_en = (top_62_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1444_in = par_reset32_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1444_write_en = (top_63_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1445_in = par_reset32_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1445_write_en = (top_64_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1446_in = par_reset32_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1446_write_en = (top_65_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1447_in = par_reset32_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1447_write_en = (top_66_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1448_in = par_reset32_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1448_write_en = (top_67_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1449_in = par_reset32_out ? 1'd0 : (top_71_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1449_write_en = (top_71_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1450_in = par_reset32_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1450_write_en = (top_72_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1451_in = par_reset32_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1451_write_en = (top_73_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1452_in = par_reset32_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1452_write_en = (top_74_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1453_in = par_reset32_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1453_write_en = (top_75_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1454_in = par_reset32_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1454_write_en = (top_76_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1455_in = par_reset32_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1455_write_en = (top_77_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1456_in = par_reset32_out ? 1'd0 : (left_17_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1456_write_en = (left_17_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1457_in = par_reset32_out ? 1'd0 : (left_26_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1457_write_en = (left_26_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1458_in = par_reset32_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1458_write_en = (left_27_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1459_in = par_reset32_out ? 1'd0 : (left_35_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1459_write_en = (left_35_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1460_in = par_reset32_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1460_write_en = (left_36_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1461_in = par_reset32_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1461_write_en = (left_37_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1462_in = par_reset32_out ? 1'd0 : (left_44_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1462_write_en = (left_44_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1463_in = par_reset32_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1463_write_en = (left_45_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1464_in = par_reset32_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1464_write_en = (left_46_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1465_in = par_reset32_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1465_write_en = (left_47_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1466_in = par_reset32_out ? 1'd0 : (left_53_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1466_write_en = (left_53_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1467_in = par_reset32_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1467_write_en = (left_54_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1468_in = par_reset32_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1468_write_en = (left_55_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1469_in = par_reset32_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1469_write_en = (left_56_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1470_in = par_reset32_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1470_write_en = (left_57_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1471_in = par_reset32_out ? 1'd0 : (left_62_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1471_write_en = (left_62_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1472_in = par_reset32_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1472_write_en = (left_63_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1473_in = par_reset32_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1473_write_en = (left_64_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1474_in = par_reset32_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1474_write_en = (left_65_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1475_in = par_reset32_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1475_write_en = (left_66_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1476_in = par_reset32_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1476_write_en = (left_67_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1477_in = par_reset32_out ? 1'd0 : (left_71_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1477_write_en = (left_71_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1478_in = par_reset32_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1478_write_en = (left_72_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1479_in = par_reset32_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1479_write_en = (left_73_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1480_in = par_reset32_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1480_write_en = (left_74_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1481_in = par_reset32_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1481_write_en = (left_75_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1482_in = par_reset32_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1482_write_en = (left_76_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_done_reg1483_in = par_reset32_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd32 & !par_reset32_out & go) ? 1'd1 : '0;
  assign par_done_reg1483_write_en = (left_77_read_done & fsm0_out == 32'd32 & !par_reset32_out & go | par_reset32_out) ? 1'd1 : '0;
  assign par_reset33_in = par_reset33_out ? 1'd0 : (par_done_reg1484_out & par_done_reg1485_out & par_done_reg1486_out & par_done_reg1487_out & par_done_reg1488_out & par_done_reg1489_out & par_done_reg1490_out & par_done_reg1491_out & par_done_reg1492_out & par_done_reg1493_out & par_done_reg1494_out & par_done_reg1495_out & par_done_reg1496_out & par_done_reg1497_out & par_done_reg1498_out & par_done_reg1499_out & par_done_reg1500_out & par_done_reg1501_out & par_done_reg1502_out & par_done_reg1503_out & par_done_reg1504_out & par_done_reg1505_out & par_done_reg1506_out & par_done_reg1507_out & par_done_reg1508_out & par_done_reg1509_out & par_done_reg1510_out & par_done_reg1511_out & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_reset33_write_en = (par_done_reg1484_out & par_done_reg1485_out & par_done_reg1486_out & par_done_reg1487_out & par_done_reg1488_out & par_done_reg1489_out & par_done_reg1490_out & par_done_reg1491_out & par_done_reg1492_out & par_done_reg1493_out & par_done_reg1494_out & par_done_reg1495_out & par_done_reg1496_out & par_done_reg1497_out & par_done_reg1498_out & par_done_reg1499_out & par_done_reg1500_out & par_done_reg1501_out & par_done_reg1502_out & par_done_reg1503_out & par_done_reg1504_out & par_done_reg1505_out & par_done_reg1506_out & par_done_reg1507_out & par_done_reg1508_out & par_done_reg1509_out & par_done_reg1510_out & par_done_reg1511_out & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1484_in = par_reset33_out ? 1'd0 : (down_17_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1484_write_en = (down_17_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1485_in = par_reset33_out ? 1'd0 : (right_26_write_done & down_26_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1485_write_en = (right_26_write_done & down_26_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1486_in = par_reset33_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1486_write_en = (down_27_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1487_in = par_reset33_out ? 1'd0 : (right_35_write_done & down_35_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1487_write_en = (right_35_write_done & down_35_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1488_in = par_reset33_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1488_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1489_in = par_reset33_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1489_write_en = (down_37_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1490_in = par_reset33_out ? 1'd0 : (right_44_write_done & down_44_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1490_write_en = (right_44_write_done & down_44_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1491_in = par_reset33_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1491_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1492_in = par_reset33_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1492_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1493_in = par_reset33_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1493_write_en = (down_47_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1494_in = par_reset33_out ? 1'd0 : (right_53_write_done & down_53_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1494_write_en = (right_53_write_done & down_53_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1495_in = par_reset33_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1495_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1496_in = par_reset33_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1496_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1497_in = par_reset33_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1497_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1498_in = par_reset33_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1498_write_en = (down_57_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1499_in = par_reset33_out ? 1'd0 : (right_62_write_done & down_62_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1499_write_en = (right_62_write_done & down_62_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1500_in = par_reset33_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1500_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1501_in = par_reset33_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1501_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1502_in = par_reset33_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1502_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1503_in = par_reset33_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1503_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1504_in = par_reset33_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1504_write_en = (down_67_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1505_in = par_reset33_out ? 1'd0 : (right_71_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1505_write_en = (right_71_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1506_in = par_reset33_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1506_write_en = (right_72_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1507_in = par_reset33_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1507_write_en = (right_73_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1508_in = par_reset33_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1508_write_en = (right_74_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1509_in = par_reset33_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1509_write_en = (right_75_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1510_in = par_reset33_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1510_write_en = (right_76_write_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_done_reg1511_in = par_reset33_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd33 & !par_reset33_out & go) ? 1'd1 : '0;
  assign par_done_reg1511_write_en = (pe_77_done & fsm0_out == 32'd33 & !par_reset33_out & go | par_reset33_out) ? 1'd1 : '0;
  assign par_reset34_in = par_reset34_out ? 1'd0 : (par_done_reg1512_out & par_done_reg1513_out & par_done_reg1514_out & par_done_reg1515_out & par_done_reg1516_out & par_done_reg1517_out & par_done_reg1518_out & par_done_reg1519_out & par_done_reg1520_out & par_done_reg1521_out & par_done_reg1522_out & par_done_reg1523_out & par_done_reg1524_out & par_done_reg1525_out & par_done_reg1526_out & par_done_reg1527_out & par_done_reg1528_out & par_done_reg1529_out & par_done_reg1530_out & par_done_reg1531_out & par_done_reg1532_out & par_done_reg1533_out & par_done_reg1534_out & par_done_reg1535_out & par_done_reg1536_out & par_done_reg1537_out & par_done_reg1538_out & par_done_reg1539_out & par_done_reg1540_out & par_done_reg1541_out & par_done_reg1542_out & par_done_reg1543_out & par_done_reg1544_out & par_done_reg1545_out & par_done_reg1546_out & par_done_reg1547_out & par_done_reg1548_out & par_done_reg1549_out & par_done_reg1550_out & par_done_reg1551_out & par_done_reg1552_out & par_done_reg1553_out & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_reset34_write_en = (par_done_reg1512_out & par_done_reg1513_out & par_done_reg1514_out & par_done_reg1515_out & par_done_reg1516_out & par_done_reg1517_out & par_done_reg1518_out & par_done_reg1519_out & par_done_reg1520_out & par_done_reg1521_out & par_done_reg1522_out & par_done_reg1523_out & par_done_reg1524_out & par_done_reg1525_out & par_done_reg1526_out & par_done_reg1527_out & par_done_reg1528_out & par_done_reg1529_out & par_done_reg1530_out & par_done_reg1531_out & par_done_reg1532_out & par_done_reg1533_out & par_done_reg1534_out & par_done_reg1535_out & par_done_reg1536_out & par_done_reg1537_out & par_done_reg1538_out & par_done_reg1539_out & par_done_reg1540_out & par_done_reg1541_out & par_done_reg1542_out & par_done_reg1543_out & par_done_reg1544_out & par_done_reg1545_out & par_done_reg1546_out & par_done_reg1547_out & par_done_reg1548_out & par_done_reg1549_out & par_done_reg1550_out & par_done_reg1551_out & par_done_reg1552_out & par_done_reg1553_out & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1512_in = par_reset34_out ? 1'd0 : (top_27_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1512_write_en = (top_27_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1513_in = par_reset34_out ? 1'd0 : (top_36_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1513_write_en = (top_36_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1514_in = par_reset34_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1514_write_en = (top_37_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1515_in = par_reset34_out ? 1'd0 : (top_45_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1515_write_en = (top_45_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1516_in = par_reset34_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1516_write_en = (top_46_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1517_in = par_reset34_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1517_write_en = (top_47_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1518_in = par_reset34_out ? 1'd0 : (top_54_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1518_write_en = (top_54_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1519_in = par_reset34_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1519_write_en = (top_55_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1520_in = par_reset34_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1520_write_en = (top_56_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1521_in = par_reset34_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1521_write_en = (top_57_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1522_in = par_reset34_out ? 1'd0 : (top_63_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1522_write_en = (top_63_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1523_in = par_reset34_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1523_write_en = (top_64_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1524_in = par_reset34_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1524_write_en = (top_65_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1525_in = par_reset34_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1525_write_en = (top_66_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1526_in = par_reset34_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1526_write_en = (top_67_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1527_in = par_reset34_out ? 1'd0 : (top_72_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1527_write_en = (top_72_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1528_in = par_reset34_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1528_write_en = (top_73_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1529_in = par_reset34_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1529_write_en = (top_74_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1530_in = par_reset34_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1530_write_en = (top_75_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1531_in = par_reset34_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1531_write_en = (top_76_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1532_in = par_reset34_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1532_write_en = (top_77_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1533_in = par_reset34_out ? 1'd0 : (left_27_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1533_write_en = (left_27_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1534_in = par_reset34_out ? 1'd0 : (left_36_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1534_write_en = (left_36_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1535_in = par_reset34_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1535_write_en = (left_37_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1536_in = par_reset34_out ? 1'd0 : (left_45_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1536_write_en = (left_45_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1537_in = par_reset34_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1537_write_en = (left_46_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1538_in = par_reset34_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1538_write_en = (left_47_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1539_in = par_reset34_out ? 1'd0 : (left_54_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1539_write_en = (left_54_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1540_in = par_reset34_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1540_write_en = (left_55_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1541_in = par_reset34_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1541_write_en = (left_56_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1542_in = par_reset34_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1542_write_en = (left_57_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1543_in = par_reset34_out ? 1'd0 : (left_63_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1543_write_en = (left_63_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1544_in = par_reset34_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1544_write_en = (left_64_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1545_in = par_reset34_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1545_write_en = (left_65_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1546_in = par_reset34_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1546_write_en = (left_66_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1547_in = par_reset34_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1547_write_en = (left_67_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1548_in = par_reset34_out ? 1'd0 : (left_72_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1548_write_en = (left_72_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1549_in = par_reset34_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1549_write_en = (left_73_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1550_in = par_reset34_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1550_write_en = (left_74_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1551_in = par_reset34_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1551_write_en = (left_75_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1552_in = par_reset34_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1552_write_en = (left_76_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_done_reg1553_in = par_reset34_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd34 & !par_reset34_out & go) ? 1'd1 : '0;
  assign par_done_reg1553_write_en = (left_77_read_done & fsm0_out == 32'd34 & !par_reset34_out & go | par_reset34_out) ? 1'd1 : '0;
  assign par_reset35_in = par_reset35_out ? 1'd0 : (par_done_reg1554_out & par_done_reg1555_out & par_done_reg1556_out & par_done_reg1557_out & par_done_reg1558_out & par_done_reg1559_out & par_done_reg1560_out & par_done_reg1561_out & par_done_reg1562_out & par_done_reg1563_out & par_done_reg1564_out & par_done_reg1565_out & par_done_reg1566_out & par_done_reg1567_out & par_done_reg1568_out & par_done_reg1569_out & par_done_reg1570_out & par_done_reg1571_out & par_done_reg1572_out & par_done_reg1573_out & par_done_reg1574_out & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_reset35_write_en = (par_done_reg1554_out & par_done_reg1555_out & par_done_reg1556_out & par_done_reg1557_out & par_done_reg1558_out & par_done_reg1559_out & par_done_reg1560_out & par_done_reg1561_out & par_done_reg1562_out & par_done_reg1563_out & par_done_reg1564_out & par_done_reg1565_out & par_done_reg1566_out & par_done_reg1567_out & par_done_reg1568_out & par_done_reg1569_out & par_done_reg1570_out & par_done_reg1571_out & par_done_reg1572_out & par_done_reg1573_out & par_done_reg1574_out & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1554_in = par_reset35_out ? 1'd0 : (down_27_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1554_write_en = (down_27_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1555_in = par_reset35_out ? 1'd0 : (right_36_write_done & down_36_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1555_write_en = (right_36_write_done & down_36_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1556_in = par_reset35_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1556_write_en = (down_37_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1557_in = par_reset35_out ? 1'd0 : (right_45_write_done & down_45_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1557_write_en = (right_45_write_done & down_45_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1558_in = par_reset35_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1558_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1559_in = par_reset35_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1559_write_en = (down_47_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1560_in = par_reset35_out ? 1'd0 : (right_54_write_done & down_54_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1560_write_en = (right_54_write_done & down_54_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1561_in = par_reset35_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1561_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1562_in = par_reset35_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1562_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1563_in = par_reset35_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1563_write_en = (down_57_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1564_in = par_reset35_out ? 1'd0 : (right_63_write_done & down_63_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1564_write_en = (right_63_write_done & down_63_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1565_in = par_reset35_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1565_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1566_in = par_reset35_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1566_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1567_in = par_reset35_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1567_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1568_in = par_reset35_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1568_write_en = (down_67_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1569_in = par_reset35_out ? 1'd0 : (right_72_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1569_write_en = (right_72_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1570_in = par_reset35_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1570_write_en = (right_73_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1571_in = par_reset35_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1571_write_en = (right_74_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1572_in = par_reset35_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1572_write_en = (right_75_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1573_in = par_reset35_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1573_write_en = (right_76_write_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_done_reg1574_in = par_reset35_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd35 & !par_reset35_out & go) ? 1'd1 : '0;
  assign par_done_reg1574_write_en = (pe_77_done & fsm0_out == 32'd35 & !par_reset35_out & go | par_reset35_out) ? 1'd1 : '0;
  assign par_reset36_in = par_reset36_out ? 1'd0 : (par_done_reg1575_out & par_done_reg1576_out & par_done_reg1577_out & par_done_reg1578_out & par_done_reg1579_out & par_done_reg1580_out & par_done_reg1581_out & par_done_reg1582_out & par_done_reg1583_out & par_done_reg1584_out & par_done_reg1585_out & par_done_reg1586_out & par_done_reg1587_out & par_done_reg1588_out & par_done_reg1589_out & par_done_reg1590_out & par_done_reg1591_out & par_done_reg1592_out & par_done_reg1593_out & par_done_reg1594_out & par_done_reg1595_out & par_done_reg1596_out & par_done_reg1597_out & par_done_reg1598_out & par_done_reg1599_out & par_done_reg1600_out & par_done_reg1601_out & par_done_reg1602_out & par_done_reg1603_out & par_done_reg1604_out & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_reset36_write_en = (par_done_reg1575_out & par_done_reg1576_out & par_done_reg1577_out & par_done_reg1578_out & par_done_reg1579_out & par_done_reg1580_out & par_done_reg1581_out & par_done_reg1582_out & par_done_reg1583_out & par_done_reg1584_out & par_done_reg1585_out & par_done_reg1586_out & par_done_reg1587_out & par_done_reg1588_out & par_done_reg1589_out & par_done_reg1590_out & par_done_reg1591_out & par_done_reg1592_out & par_done_reg1593_out & par_done_reg1594_out & par_done_reg1595_out & par_done_reg1596_out & par_done_reg1597_out & par_done_reg1598_out & par_done_reg1599_out & par_done_reg1600_out & par_done_reg1601_out & par_done_reg1602_out & par_done_reg1603_out & par_done_reg1604_out & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1575_in = par_reset36_out ? 1'd0 : (top_37_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1575_write_en = (top_37_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1576_in = par_reset36_out ? 1'd0 : (top_46_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1576_write_en = (top_46_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1577_in = par_reset36_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1577_write_en = (top_47_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1578_in = par_reset36_out ? 1'd0 : (top_55_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1578_write_en = (top_55_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1579_in = par_reset36_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1579_write_en = (top_56_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1580_in = par_reset36_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1580_write_en = (top_57_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1581_in = par_reset36_out ? 1'd0 : (top_64_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1581_write_en = (top_64_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1582_in = par_reset36_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1582_write_en = (top_65_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1583_in = par_reset36_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1583_write_en = (top_66_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1584_in = par_reset36_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1584_write_en = (top_67_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1585_in = par_reset36_out ? 1'd0 : (top_73_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1585_write_en = (top_73_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1586_in = par_reset36_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1586_write_en = (top_74_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1587_in = par_reset36_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1587_write_en = (top_75_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1588_in = par_reset36_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1588_write_en = (top_76_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1589_in = par_reset36_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1589_write_en = (top_77_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1590_in = par_reset36_out ? 1'd0 : (left_37_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1590_write_en = (left_37_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1591_in = par_reset36_out ? 1'd0 : (left_46_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1591_write_en = (left_46_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1592_in = par_reset36_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1592_write_en = (left_47_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1593_in = par_reset36_out ? 1'd0 : (left_55_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1593_write_en = (left_55_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1594_in = par_reset36_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1594_write_en = (left_56_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1595_in = par_reset36_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1595_write_en = (left_57_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1596_in = par_reset36_out ? 1'd0 : (left_64_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1596_write_en = (left_64_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1597_in = par_reset36_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1597_write_en = (left_65_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1598_in = par_reset36_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1598_write_en = (left_66_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1599_in = par_reset36_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1599_write_en = (left_67_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1600_in = par_reset36_out ? 1'd0 : (left_73_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1600_write_en = (left_73_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1601_in = par_reset36_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1601_write_en = (left_74_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1602_in = par_reset36_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1602_write_en = (left_75_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1603_in = par_reset36_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1603_write_en = (left_76_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_done_reg1604_in = par_reset36_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd36 & !par_reset36_out & go) ? 1'd1 : '0;
  assign par_done_reg1604_write_en = (left_77_read_done & fsm0_out == 32'd36 & !par_reset36_out & go | par_reset36_out) ? 1'd1 : '0;
  assign par_reset37_in = par_reset37_out ? 1'd0 : (par_done_reg1605_out & par_done_reg1606_out & par_done_reg1607_out & par_done_reg1608_out & par_done_reg1609_out & par_done_reg1610_out & par_done_reg1611_out & par_done_reg1612_out & par_done_reg1613_out & par_done_reg1614_out & par_done_reg1615_out & par_done_reg1616_out & par_done_reg1617_out & par_done_reg1618_out & par_done_reg1619_out & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_reset37_write_en = (par_done_reg1605_out & par_done_reg1606_out & par_done_reg1607_out & par_done_reg1608_out & par_done_reg1609_out & par_done_reg1610_out & par_done_reg1611_out & par_done_reg1612_out & par_done_reg1613_out & par_done_reg1614_out & par_done_reg1615_out & par_done_reg1616_out & par_done_reg1617_out & par_done_reg1618_out & par_done_reg1619_out & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1605_in = par_reset37_out ? 1'd0 : (down_37_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1605_write_en = (down_37_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1606_in = par_reset37_out ? 1'd0 : (right_46_write_done & down_46_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1606_write_en = (right_46_write_done & down_46_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1607_in = par_reset37_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1607_write_en = (down_47_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1608_in = par_reset37_out ? 1'd0 : (right_55_write_done & down_55_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1608_write_en = (right_55_write_done & down_55_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1609_in = par_reset37_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1609_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1610_in = par_reset37_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1610_write_en = (down_57_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1611_in = par_reset37_out ? 1'd0 : (right_64_write_done & down_64_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1611_write_en = (right_64_write_done & down_64_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1612_in = par_reset37_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1612_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1613_in = par_reset37_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1613_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1614_in = par_reset37_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1614_write_en = (down_67_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1615_in = par_reset37_out ? 1'd0 : (right_73_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1615_write_en = (right_73_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1616_in = par_reset37_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1616_write_en = (right_74_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1617_in = par_reset37_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1617_write_en = (right_75_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1618_in = par_reset37_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1618_write_en = (right_76_write_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_done_reg1619_in = par_reset37_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd37 & !par_reset37_out & go) ? 1'd1 : '0;
  assign par_done_reg1619_write_en = (pe_77_done & fsm0_out == 32'd37 & !par_reset37_out & go | par_reset37_out) ? 1'd1 : '0;
  assign par_reset38_in = par_reset38_out ? 1'd0 : (par_done_reg1620_out & par_done_reg1621_out & par_done_reg1622_out & par_done_reg1623_out & par_done_reg1624_out & par_done_reg1625_out & par_done_reg1626_out & par_done_reg1627_out & par_done_reg1628_out & par_done_reg1629_out & par_done_reg1630_out & par_done_reg1631_out & par_done_reg1632_out & par_done_reg1633_out & par_done_reg1634_out & par_done_reg1635_out & par_done_reg1636_out & par_done_reg1637_out & par_done_reg1638_out & par_done_reg1639_out & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_reset38_write_en = (par_done_reg1620_out & par_done_reg1621_out & par_done_reg1622_out & par_done_reg1623_out & par_done_reg1624_out & par_done_reg1625_out & par_done_reg1626_out & par_done_reg1627_out & par_done_reg1628_out & par_done_reg1629_out & par_done_reg1630_out & par_done_reg1631_out & par_done_reg1632_out & par_done_reg1633_out & par_done_reg1634_out & par_done_reg1635_out & par_done_reg1636_out & par_done_reg1637_out & par_done_reg1638_out & par_done_reg1639_out & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1620_in = par_reset38_out ? 1'd0 : (top_47_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1620_write_en = (top_47_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1621_in = par_reset38_out ? 1'd0 : (top_56_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1621_write_en = (top_56_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1622_in = par_reset38_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1622_write_en = (top_57_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1623_in = par_reset38_out ? 1'd0 : (top_65_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1623_write_en = (top_65_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1624_in = par_reset38_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1624_write_en = (top_66_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1625_in = par_reset38_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1625_write_en = (top_67_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1626_in = par_reset38_out ? 1'd0 : (top_74_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1626_write_en = (top_74_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1627_in = par_reset38_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1627_write_en = (top_75_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1628_in = par_reset38_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1628_write_en = (top_76_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1629_in = par_reset38_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1629_write_en = (top_77_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1630_in = par_reset38_out ? 1'd0 : (left_47_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1630_write_en = (left_47_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1631_in = par_reset38_out ? 1'd0 : (left_56_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1631_write_en = (left_56_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1632_in = par_reset38_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1632_write_en = (left_57_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1633_in = par_reset38_out ? 1'd0 : (left_65_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1633_write_en = (left_65_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1634_in = par_reset38_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1634_write_en = (left_66_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1635_in = par_reset38_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1635_write_en = (left_67_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1636_in = par_reset38_out ? 1'd0 : (left_74_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1636_write_en = (left_74_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1637_in = par_reset38_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1637_write_en = (left_75_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1638_in = par_reset38_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1638_write_en = (left_76_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_done_reg1639_in = par_reset38_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd38 & !par_reset38_out & go) ? 1'd1 : '0;
  assign par_done_reg1639_write_en = (left_77_read_done & fsm0_out == 32'd38 & !par_reset38_out & go | par_reset38_out) ? 1'd1 : '0;
  assign par_reset39_in = par_reset39_out ? 1'd0 : (par_done_reg1640_out & par_done_reg1641_out & par_done_reg1642_out & par_done_reg1643_out & par_done_reg1644_out & par_done_reg1645_out & par_done_reg1646_out & par_done_reg1647_out & par_done_reg1648_out & par_done_reg1649_out & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_reset39_write_en = (par_done_reg1640_out & par_done_reg1641_out & par_done_reg1642_out & par_done_reg1643_out & par_done_reg1644_out & par_done_reg1645_out & par_done_reg1646_out & par_done_reg1647_out & par_done_reg1648_out & par_done_reg1649_out & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1640_in = par_reset39_out ? 1'd0 : (down_47_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1640_write_en = (down_47_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1641_in = par_reset39_out ? 1'd0 : (right_56_write_done & down_56_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1641_write_en = (right_56_write_done & down_56_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1642_in = par_reset39_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1642_write_en = (down_57_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1643_in = par_reset39_out ? 1'd0 : (right_65_write_done & down_65_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1643_write_en = (right_65_write_done & down_65_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1644_in = par_reset39_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1644_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1645_in = par_reset39_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1645_write_en = (down_67_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1646_in = par_reset39_out ? 1'd0 : (right_74_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1646_write_en = (right_74_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1647_in = par_reset39_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1647_write_en = (right_75_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1648_in = par_reset39_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1648_write_en = (right_76_write_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_done_reg1649_in = par_reset39_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd39 & !par_reset39_out & go) ? 1'd1 : '0;
  assign par_done_reg1649_write_en = (pe_77_done & fsm0_out == 32'd39 & !par_reset39_out & go | par_reset39_out) ? 1'd1 : '0;
  assign par_reset40_in = par_reset40_out ? 1'd0 : (par_done_reg1650_out & par_done_reg1651_out & par_done_reg1652_out & par_done_reg1653_out & par_done_reg1654_out & par_done_reg1655_out & par_done_reg1656_out & par_done_reg1657_out & par_done_reg1658_out & par_done_reg1659_out & par_done_reg1660_out & par_done_reg1661_out & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_reset40_write_en = (par_done_reg1650_out & par_done_reg1651_out & par_done_reg1652_out & par_done_reg1653_out & par_done_reg1654_out & par_done_reg1655_out & par_done_reg1656_out & par_done_reg1657_out & par_done_reg1658_out & par_done_reg1659_out & par_done_reg1660_out & par_done_reg1661_out & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1650_in = par_reset40_out ? 1'd0 : (top_57_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1650_write_en = (top_57_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1651_in = par_reset40_out ? 1'd0 : (top_66_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1651_write_en = (top_66_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1652_in = par_reset40_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1652_write_en = (top_67_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1653_in = par_reset40_out ? 1'd0 : (top_75_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1653_write_en = (top_75_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1654_in = par_reset40_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1654_write_en = (top_76_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1655_in = par_reset40_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1655_write_en = (top_77_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1656_in = par_reset40_out ? 1'd0 : (left_57_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1656_write_en = (left_57_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1657_in = par_reset40_out ? 1'd0 : (left_66_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1657_write_en = (left_66_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1658_in = par_reset40_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1658_write_en = (left_67_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1659_in = par_reset40_out ? 1'd0 : (left_75_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1659_write_en = (left_75_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1660_in = par_reset40_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1660_write_en = (left_76_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_done_reg1661_in = par_reset40_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd40 & !par_reset40_out & go) ? 1'd1 : '0;
  assign par_done_reg1661_write_en = (left_77_read_done & fsm0_out == 32'd40 & !par_reset40_out & go | par_reset40_out) ? 1'd1 : '0;
  assign par_reset41_in = par_reset41_out ? 1'd0 : (par_done_reg1662_out & par_done_reg1663_out & par_done_reg1664_out & par_done_reg1665_out & par_done_reg1666_out & par_done_reg1667_out & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_reset41_write_en = (par_done_reg1662_out & par_done_reg1663_out & par_done_reg1664_out & par_done_reg1665_out & par_done_reg1666_out & par_done_reg1667_out & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_done_reg1662_in = par_reset41_out ? 1'd0 : (down_57_write_done & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_done_reg1662_write_en = (down_57_write_done & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_done_reg1663_in = par_reset41_out ? 1'd0 : (right_66_write_done & down_66_write_done & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_done_reg1663_write_en = (right_66_write_done & down_66_write_done & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_done_reg1664_in = par_reset41_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_done_reg1664_write_en = (down_67_write_done & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_done_reg1665_in = par_reset41_out ? 1'd0 : (right_75_write_done & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_done_reg1665_write_en = (right_75_write_done & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_done_reg1666_in = par_reset41_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_done_reg1666_write_en = (right_76_write_done & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_done_reg1667_in = par_reset41_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd41 & !par_reset41_out & go) ? 1'd1 : '0;
  assign par_done_reg1667_write_en = (pe_77_done & fsm0_out == 32'd41 & !par_reset41_out & go | par_reset41_out) ? 1'd1 : '0;
  assign par_reset42_in = par_reset42_out ? 1'd0 : (par_done_reg1668_out & par_done_reg1669_out & par_done_reg1670_out & par_done_reg1671_out & par_done_reg1672_out & par_done_reg1673_out & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_reset42_write_en = (par_done_reg1668_out & par_done_reg1669_out & par_done_reg1670_out & par_done_reg1671_out & par_done_reg1672_out & par_done_reg1673_out & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_done_reg1668_in = par_reset42_out ? 1'd0 : (top_67_read_done & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_done_reg1668_write_en = (top_67_read_done & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_done_reg1669_in = par_reset42_out ? 1'd0 : (top_76_read_done & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_done_reg1669_write_en = (top_76_read_done & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_done_reg1670_in = par_reset42_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_done_reg1670_write_en = (top_77_read_done & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_done_reg1671_in = par_reset42_out ? 1'd0 : (left_67_read_done & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_done_reg1671_write_en = (left_67_read_done & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_done_reg1672_in = par_reset42_out ? 1'd0 : (left_76_read_done & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_done_reg1672_write_en = (left_76_read_done & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_done_reg1673_in = par_reset42_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd42 & !par_reset42_out & go) ? 1'd1 : '0;
  assign par_done_reg1673_write_en = (left_77_read_done & fsm0_out == 32'd42 & !par_reset42_out & go | par_reset42_out) ? 1'd1 : '0;
  assign par_reset43_in = par_reset43_out ? 1'd0 : (par_done_reg1674_out & par_done_reg1675_out & par_done_reg1676_out & fsm0_out == 32'd43 & !par_reset43_out & go) ? 1'd1 : '0;
  assign par_reset43_write_en = (par_done_reg1674_out & par_done_reg1675_out & par_done_reg1676_out & fsm0_out == 32'd43 & !par_reset43_out & go | par_reset43_out) ? 1'd1 : '0;
  assign par_done_reg1674_in = par_reset43_out ? 1'd0 : (down_67_write_done & fsm0_out == 32'd43 & !par_reset43_out & go) ? 1'd1 : '0;
  assign par_done_reg1674_write_en = (down_67_write_done & fsm0_out == 32'd43 & !par_reset43_out & go | par_reset43_out) ? 1'd1 : '0;
  assign par_done_reg1675_in = par_reset43_out ? 1'd0 : (right_76_write_done & fsm0_out == 32'd43 & !par_reset43_out & go) ? 1'd1 : '0;
  assign par_done_reg1675_write_en = (right_76_write_done & fsm0_out == 32'd43 & !par_reset43_out & go | par_reset43_out) ? 1'd1 : '0;
  assign par_done_reg1676_in = par_reset43_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd43 & !par_reset43_out & go) ? 1'd1 : '0;
  assign par_done_reg1676_write_en = (pe_77_done & fsm0_out == 32'd43 & !par_reset43_out & go | par_reset43_out) ? 1'd1 : '0;
  assign par_reset44_in = par_reset44_out ? 1'd0 : (par_done_reg1677_out & par_done_reg1678_out & fsm0_out == 32'd44 & !par_reset44_out & go) ? 1'd1 : '0;
  assign par_reset44_write_en = (par_done_reg1677_out & par_done_reg1678_out & fsm0_out == 32'd44 & !par_reset44_out & go | par_reset44_out) ? 1'd1 : '0;
  assign par_done_reg1677_in = par_reset44_out ? 1'd0 : (top_77_read_done & fsm0_out == 32'd44 & !par_reset44_out & go) ? 1'd1 : '0;
  assign par_done_reg1677_write_en = (top_77_read_done & fsm0_out == 32'd44 & !par_reset44_out & go | par_reset44_out) ? 1'd1 : '0;
  assign par_done_reg1678_in = par_reset44_out ? 1'd0 : (left_77_read_done & fsm0_out == 32'd44 & !par_reset44_out & go) ? 1'd1 : '0;
  assign par_done_reg1678_write_en = (left_77_read_done & fsm0_out == 32'd44 & !par_reset44_out & go | par_reset44_out) ? 1'd1 : '0;
  assign par_reset45_in = par_reset45_out ? 1'd0 : (par_done_reg1679_out & fsm0_out == 32'd45 & !par_reset45_out & go) ? 1'd1 : '0;
  assign par_reset45_write_en = (par_done_reg1679_out & fsm0_out == 32'd45 & !par_reset45_out & go | par_reset45_out) ? 1'd1 : '0;
  assign par_done_reg1679_in = par_reset45_out ? 1'd0 : (pe_77_done & fsm0_out == 32'd45 & !par_reset45_out & go) ? 1'd1 : '0;
  assign par_done_reg1679_write_en = (pe_77_done & fsm0_out == 32'd45 & !par_reset45_out & go | par_reset45_out) ? 1'd1 : '0;
  assign fsm0_in = (fsm0_out == 32'd87 & out_mem_done & go) ? 32'd88 : (fsm0_out == 32'd86 & out_mem_done & go) ? 32'd87 : (fsm0_out == 32'd85 & out_mem_done & go) ? 32'd86 : (fsm0_out == 32'd84 & out_mem_done & go) ? 32'd85 : (fsm0_out == 32'd83 & out_mem_done & go) ? 32'd84 : (fsm0_out == 32'd82 & out_mem_done & go) ? 32'd83 : (fsm0_out == 32'd81 & out_mem_done & go) ? 32'd82 : (fsm0_out == 32'd80 & out_mem_done & go) ? 32'd81 : (fsm0_out == 32'd79 & out_mem_done & go) ? 32'd80 : (fsm0_out == 32'd78 & out_mem_done & go) ? 32'd79 : (fsm0_out == 32'd77 & out_mem_done & go) ? 32'd78 : (fsm0_out == 32'd76 & out_mem_done & go) ? 32'd77 : (fsm0_out == 32'd75 & out_mem_done & go) ? 32'd76 : (fsm0_out == 32'd74 & out_mem_done & go) ? 32'd75 : (fsm0_out == 32'd73 & out_mem_done & go) ? 32'd74 : (fsm0_out == 32'd72 & out_mem_done & go) ? 32'd73 : (fsm0_out == 32'd71 & out_mem_done & go) ? 32'd72 : (fsm0_out == 32'd70 & out_mem_done & go) ? 32'd71 : (fsm0_out == 32'd69 & out_mem_done & go) ? 32'd70 : (fsm0_out == 32'd68 & out_mem_done & go) ? 32'd69 : (fsm0_out == 32'd67 & out_mem_done & go) ? 32'd68 : (fsm0_out == 32'd66 & out_mem_done & go) ? 32'd67 : (fsm0_out == 32'd65 & out_mem_done & go) ? 32'd66 : (fsm0_out == 32'd64 & out_mem_done & go) ? 32'd65 : (fsm0_out == 32'd63 & out_mem_done & go) ? 32'd64 : (fsm0_out == 32'd62 & out_mem_done & go) ? 32'd63 : (fsm0_out == 32'd61 & out_mem_done & go) ? 32'd62 : (fsm0_out == 32'd60 & out_mem_done & go) ? 32'd61 : (fsm0_out == 32'd59 & out_mem_done & go) ? 32'd60 : (fsm0_out == 32'd58 & out_mem_done & go) ? 32'd59 : (fsm0_out == 32'd57 & out_mem_done & go) ? 32'd58 : (fsm0_out == 32'd56 & out_mem_done & go) ? 32'd57 : (fsm0_out == 32'd55 & out_mem_done & go) ? 32'd56 : (fsm0_out == 32'd54 & out_mem_done & go) ? 32'd55 : (fsm0_out == 32'd53 & out_mem_done & go) ? 32'd54 : (fsm0_out == 32'd52 & out_mem_done & go) ? 32'd53 : (fsm0_out == 32'd51 & out_mem_done & go) ? 32'd52 : (fsm0_out == 32'd50 & out_mem_done & go) ? 32'd51 : (fsm0_out == 32'd49 & out_mem_done & go) ? 32'd50 : (fsm0_out == 32'd48 & out_mem_done & go) ? 32'd49 : (fsm0_out == 32'd47 & out_mem_done & go) ? 32'd48 : (fsm0_out == 32'd46 & out_mem_done & go) ? 32'd47 : (fsm0_out == 32'd45 & par_reset45_out & go) ? 32'd46 : (fsm0_out == 32'd44 & par_reset44_out & go) ? 32'd45 : (fsm0_out == 32'd43 & par_reset43_out & go) ? 32'd44 : (fsm0_out == 32'd42 & par_reset42_out & go) ? 32'd43 : (fsm0_out == 32'd41 & par_reset41_out & go) ? 32'd42 : (fsm0_out == 32'd40 & par_reset40_out & go) ? 32'd41 : (fsm0_out == 32'd39 & par_reset39_out & go) ? 32'd40 : (fsm0_out == 32'd38 & par_reset38_out & go) ? 32'd39 : (fsm0_out == 32'd37 & par_reset37_out & go) ? 32'd38 : (fsm0_out == 32'd36 & par_reset36_out & go) ? 32'd37 : (fsm0_out == 32'd35 & par_reset35_out & go) ? 32'd36 : (fsm0_out == 32'd34 & par_reset34_out & go) ? 32'd35 : (fsm0_out == 32'd33 & par_reset33_out & go) ? 32'd34 : (fsm0_out == 32'd32 & par_reset32_out & go) ? 32'd33 : (fsm0_out == 32'd31 & par_reset31_out & go) ? 32'd32 : (fsm0_out == 32'd30 & par_reset30_out & go) ? 32'd31 : (fsm0_out == 32'd29 & par_reset29_out & go) ? 32'd30 : (fsm0_out == 32'd28 & par_reset28_out & go) ? 32'd29 : (fsm0_out == 32'd27 & par_reset27_out & go) ? 32'd28 : (fsm0_out == 32'd26 & par_reset26_out & go) ? 32'd27 : (fsm0_out == 32'd25 & par_reset25_out & go) ? 32'd26 : (fsm0_out == 32'd24 & par_reset24_out & go) ? 32'd25 : (fsm0_out == 32'd23 & par_reset23_out & go) ? 32'd24 : (fsm0_out == 32'd22 & par_reset22_out & go) ? 32'd23 : (fsm0_out == 32'd21 & par_reset21_out & go) ? 32'd22 : (fsm0_out == 32'd20 & par_reset20_out & go) ? 32'd21 : (fsm0_out == 32'd19 & par_reset19_out & go) ? 32'd20 : (fsm0_out == 32'd18 & par_reset18_out & go) ? 32'd19 : (fsm0_out == 32'd17 & par_reset17_out & go) ? 32'd18 : (fsm0_out == 32'd16 & par_reset16_out & go) ? 32'd17 : (fsm0_out == 32'd15 & par_reset15_out & go) ? 32'd16 : (fsm0_out == 32'd14 & par_reset14_out & go) ? 32'd15 : (fsm0_out == 32'd13 & par_reset13_out & go) ? 32'd14 : (fsm0_out == 32'd12 & par_reset12_out & go) ? 32'd13 : (fsm0_out == 32'd11 & par_reset11_out & go) ? 32'd12 : (fsm0_out == 32'd10 & par_reset10_out & go) ? 32'd11 : (fsm0_out == 32'd9 & par_reset9_out & go) ? 32'd10 : (fsm0_out == 32'd8 & par_reset8_out & go) ? 32'd9 : (fsm0_out == 32'd7 & par_reset7_out & go) ? 32'd8 : (fsm0_out == 32'd6 & par_reset6_out & go) ? 32'd7 : (fsm0_out == 32'd5 & par_reset5_out & go) ? 32'd6 : (fsm0_out == 32'd4 & par_reset4_out & go) ? 32'd5 : (fsm0_out == 32'd3 & par_reset3_out & go) ? 32'd4 : (fsm0_out == 32'd2 & par_reset2_out & go) ? 32'd3 : (fsm0_out == 32'd1 & par_reset1_out & go) ? 32'd2 : (fsm0_out == 32'd109 & out_mem_done & go) ? 32'd110 : (fsm0_out == 32'd108 & out_mem_done & go) ? 32'd109 : (fsm0_out == 32'd0 & par_reset0_out & go) ? 32'd1 : (fsm0_out == 32'd107 & out_mem_done & go) ? 32'd108 : (fsm0_out == 32'd106 & out_mem_done & go) ? 32'd107 : (fsm0_out == 32'd105 & out_mem_done & go) ? 32'd106 : (fsm0_out == 32'd104 & out_mem_done & go) ? 32'd105 : (fsm0_out == 32'd103 & out_mem_done & go) ? 32'd104 : (fsm0_out == 32'd102 & out_mem_done & go) ? 32'd103 : (fsm0_out == 32'd101 & out_mem_done & go) ? 32'd102 : (fsm0_out == 32'd100 & out_mem_done & go) ? 32'd101 : (fsm0_out == 32'd99 & out_mem_done & go) ? 32'd100 : (fsm0_out == 32'd98 & out_mem_done & go) ? 32'd99 : (fsm0_out == 32'd110) ? 32'd0 : (fsm0_out == 32'd97 & out_mem_done & go) ? 32'd98 : (fsm0_out == 32'd96 & out_mem_done & go) ? 32'd97 : (fsm0_out == 32'd95 & out_mem_done & go) ? 32'd96 : (fsm0_out == 32'd94 & out_mem_done & go) ? 32'd95 : (fsm0_out == 32'd93 & out_mem_done & go) ? 32'd94 : (fsm0_out == 32'd92 & out_mem_done & go) ? 32'd93 : (fsm0_out == 32'd91 & out_mem_done & go) ? 32'd92 : (fsm0_out == 32'd90 & out_mem_done & go) ? 32'd91 : (fsm0_out == 32'd89 & out_mem_done & go) ? 32'd90 : (fsm0_out == 32'd88 & out_mem_done & go) ? 32'd89 : '0;
  assign fsm0_write_en = (fsm0_out == 32'd0 & par_reset0_out & go | fsm0_out == 32'd1 & par_reset1_out & go | fsm0_out == 32'd2 & par_reset2_out & go | fsm0_out == 32'd3 & par_reset3_out & go | fsm0_out == 32'd4 & par_reset4_out & go | fsm0_out == 32'd5 & par_reset5_out & go | fsm0_out == 32'd6 & par_reset6_out & go | fsm0_out == 32'd7 & par_reset7_out & go | fsm0_out == 32'd8 & par_reset8_out & go | fsm0_out == 32'd9 & par_reset9_out & go | fsm0_out == 32'd10 & par_reset10_out & go | fsm0_out == 32'd11 & par_reset11_out & go | fsm0_out == 32'd12 & par_reset12_out & go | fsm0_out == 32'd13 & par_reset13_out & go | fsm0_out == 32'd14 & par_reset14_out & go | fsm0_out == 32'd15 & par_reset15_out & go | fsm0_out == 32'd16 & par_reset16_out & go | fsm0_out == 32'd17 & par_reset17_out & go | fsm0_out == 32'd18 & par_reset18_out & go | fsm0_out == 32'd19 & par_reset19_out & go | fsm0_out == 32'd20 & par_reset20_out & go | fsm0_out == 32'd21 & par_reset21_out & go | fsm0_out == 32'd22 & par_reset22_out & go | fsm0_out == 32'd23 & par_reset23_out & go | fsm0_out == 32'd24 & par_reset24_out & go | fsm0_out == 32'd25 & par_reset25_out & go | fsm0_out == 32'd26 & par_reset26_out & go | fsm0_out == 32'd27 & par_reset27_out & go | fsm0_out == 32'd28 & par_reset28_out & go | fsm0_out == 32'd29 & par_reset29_out & go | fsm0_out == 32'd30 & par_reset30_out & go | fsm0_out == 32'd31 & par_reset31_out & go | fsm0_out == 32'd32 & par_reset32_out & go | fsm0_out == 32'd33 & par_reset33_out & go | fsm0_out == 32'd34 & par_reset34_out & go | fsm0_out == 32'd35 & par_reset35_out & go | fsm0_out == 32'd36 & par_reset36_out & go | fsm0_out == 32'd37 & par_reset37_out & go | fsm0_out == 32'd38 & par_reset38_out & go | fsm0_out == 32'd39 & par_reset39_out & go | fsm0_out == 32'd40 & par_reset40_out & go | fsm0_out == 32'd41 & par_reset41_out & go | fsm0_out == 32'd42 & par_reset42_out & go | fsm0_out == 32'd43 & par_reset43_out & go | fsm0_out == 32'd44 & par_reset44_out & go | fsm0_out == 32'd45 & par_reset45_out & go | fsm0_out == 32'd46 & out_mem_done & go | fsm0_out == 32'd47 & out_mem_done & go | fsm0_out == 32'd48 & out_mem_done & go | fsm0_out == 32'd49 & out_mem_done & go | fsm0_out == 32'd50 & out_mem_done & go | fsm0_out == 32'd51 & out_mem_done & go | fsm0_out == 32'd52 & out_mem_done & go | fsm0_out == 32'd53 & out_mem_done & go | fsm0_out == 32'd54 & out_mem_done & go | fsm0_out == 32'd55 & out_mem_done & go | fsm0_out == 32'd56 & out_mem_done & go | fsm0_out == 32'd57 & out_mem_done & go | fsm0_out == 32'd58 & out_mem_done & go | fsm0_out == 32'd59 & out_mem_done & go | fsm0_out == 32'd60 & out_mem_done & go | fsm0_out == 32'd61 & out_mem_done & go | fsm0_out == 32'd62 & out_mem_done & go | fsm0_out == 32'd63 & out_mem_done & go | fsm0_out == 32'd64 & out_mem_done & go | fsm0_out == 32'd65 & out_mem_done & go | fsm0_out == 32'd66 & out_mem_done & go | fsm0_out == 32'd67 & out_mem_done & go | fsm0_out == 32'd68 & out_mem_done & go | fsm0_out == 32'd69 & out_mem_done & go | fsm0_out == 32'd70 & out_mem_done & go | fsm0_out == 32'd71 & out_mem_done & go | fsm0_out == 32'd72 & out_mem_done & go | fsm0_out == 32'd73 & out_mem_done & go | fsm0_out == 32'd74 & out_mem_done & go | fsm0_out == 32'd75 & out_mem_done & go | fsm0_out == 32'd76 & out_mem_done & go | fsm0_out == 32'd77 & out_mem_done & go | fsm0_out == 32'd78 & out_mem_done & go | fsm0_out == 32'd79 & out_mem_done & go | fsm0_out == 32'd80 & out_mem_done & go | fsm0_out == 32'd81 & out_mem_done & go | fsm0_out == 32'd82 & out_mem_done & go | fsm0_out == 32'd83 & out_mem_done & go | fsm0_out == 32'd84 & out_mem_done & go | fsm0_out == 32'd85 & out_mem_done & go | fsm0_out == 32'd86 & out_mem_done & go | fsm0_out == 32'd87 & out_mem_done & go | fsm0_out == 32'd88 & out_mem_done & go | fsm0_out == 32'd89 & out_mem_done & go | fsm0_out == 32'd90 & out_mem_done & go | fsm0_out == 32'd91 & out_mem_done & go | fsm0_out == 32'd92 & out_mem_done & go | fsm0_out == 32'd93 & out_mem_done & go | fsm0_out == 32'd94 & out_mem_done & go | fsm0_out == 32'd95 & out_mem_done & go | fsm0_out == 32'd96 & out_mem_done & go | fsm0_out == 32'd97 & out_mem_done & go | fsm0_out == 32'd98 & out_mem_done & go | fsm0_out == 32'd99 & out_mem_done & go | fsm0_out == 32'd100 & out_mem_done & go | fsm0_out == 32'd101 & out_mem_done & go | fsm0_out == 32'd102 & out_mem_done & go | fsm0_out == 32'd103 & out_mem_done & go | fsm0_out == 32'd104 & out_mem_done & go | fsm0_out == 32'd105 & out_mem_done & go | fsm0_out == 32'd106 & out_mem_done & go | fsm0_out == 32'd107 & out_mem_done & go | fsm0_out == 32'd108 & out_mem_done & go | fsm0_out == 32'd109 & out_mem_done & go | fsm0_out == 32'd110) ? 1'd1 : '0;
endmodule // end main