module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule
module std_const
  #(parameter width = 32,
    parameter value = 0)
   (output logic [width - 1:0] out);
  assign out = value;
endmodule
module std_le
  #(parameter width = 32)
  (input logic [width-1:0] left,
   input logic [width-1:0] right,
   output logic            out);
  assign out = left <= right;
endmodule
module std_mem_d1
  #(parameter width = 32,
    parameter size = 16,
    parameter idx_size = 4)
   (input logic [idx_size-1:0] addr0,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  logic [width-1:0]  mem[size-1:0];

  /* verilator lint_off WIDTH */
  assign read_data = mem[addr0];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule
module std_mem_d2
  #(parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4)
   (input logic [d0_idx_size-1:0] addr0,
    input logic [d1_idx_size-1:0] addr1,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  /* verilator lint_off WIDTH */
  logic [width-1:0]  mem[d0_size-1:0][d1_size-1:0];

  assign read_data = mem[addr0][addr1];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule
module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule
module std_rsh
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left >> right;
endmodule
module kernel (
    input logic go,
    input logic clk,
    output logic done,
    output logic [6:0] A_int0_0_addr0,
    output logic [6:0] A_int0_0_addr1,
    output logic [31:0] A_int0_0_write_data,
    output logic A_int0_0_write_en,
    output logic A_int0_0_clk,
    input logic [31:0] A_int0_0_read_data,
    input logic A_int0_0_done,
    output logic alpha_int0_addr0,
    output logic [31:0] alpha_int0_write_data,
    output logic alpha_int0_write_en,
    output logic alpha_int0_clk,
    input logic [31:0] alpha_int0_read_data,
    input logic alpha_int0_done,
    output logic beta_int0_addr0,
    output logic [31:0] beta_int0_write_data,
    output logic beta_int0_write_en,
    output logic beta_int0_clk,
    input logic [31:0] beta_int0_read_data,
    input logic beta_int0_done,
    output logic [6:0] u1_int0_addr0,
    output logic [31:0] u1_int0_write_data,
    output logic u1_int0_write_en,
    output logic u1_int0_clk,
    input logic [31:0] u1_int0_read_data,
    input logic u1_int0_done,
    output logic [6:0] u2_int0_addr0,
    output logic [31:0] u2_int0_write_data,
    output logic u2_int0_write_en,
    output logic u2_int0_clk,
    input logic [31:0] u2_int0_read_data,
    input logic u2_int0_done,
    output logic [6:0] v1_int0_addr0,
    output logic [31:0] v1_int0_write_data,
    output logic v1_int0_write_en,
    output logic v1_int0_clk,
    input logic [31:0] v1_int0_read_data,
    input logic v1_int0_done,
    output logic [6:0] v2_int0_addr0,
    output logic [31:0] v2_int0_write_data,
    output logic v2_int0_write_en,
    output logic v2_int0_clk,
    input logic [31:0] v2_int0_read_data,
    input logic v2_int0_done,
    output logic [6:0] w_int0_addr0,
    output logic [31:0] w_int0_write_data,
    output logic w_int0_write_en,
    output logic w_int0_clk,
    input logic [31:0] w_int0_read_data,
    input logic w_int0_done,
    output logic [6:0] x_int0_addr0,
    output logic [31:0] x_int0_write_data,
    output logic x_int0_write_en,
    output logic x_int0_clk,
    input logic [31:0] x_int0_read_data,
    input logic x_int0_done,
    output logic [6:0] y_int0_addr0,
    output logic [31:0] y_int0_write_data,
    output logic y_int0_write_en,
    output logic y_int0_clk,
    input logic [31:0] y_int0_read_data,
    input logic y_int0_done,
    output logic [6:0] z_int0_addr0,
    output logic [31:0] z_int0_write_data,
    output logic z_int0_write_en,
    output logic z_int0_clk,
    input logic [31:0] z_int0_read_data,
    input logic z_int0_done
);
    import "DPI-C" function string futil_getenv (input string env_var);
    string DATA;
    initial begin
        DATA = futil_getenv("DATA");
        $fdisplay(2, "DATA (path to meminit files): %s", DATA);
        $readmemh({DATA, "/A0_0.dat"}, A0_0.mem);
        $readmemh({DATA, "/u10.dat"}, u10.mem);
        $readmemh({DATA, "/u20.dat"}, u20.mem);
        $readmemh({DATA, "/v10.dat"}, v10.mem);
        $readmemh({DATA, "/v20.dat"}, v20.mem);
        $readmemh({DATA, "/w0.dat"}, w0.mem);
        $readmemh({DATA, "/x0.dat"}, x0.mem);
        $readmemh({DATA, "/y0.dat"}, y0.mem);
        $readmemh({DATA, "/z0.dat"}, z0.mem);
    end
    final begin
        $writememh({DATA, "/A0_0.out"}, A0_0.mem);
        $writememh({DATA, "/u10.out"}, u10.mem);
        $writememh({DATA, "/u20.out"}, u20.mem);
        $writememh({DATA, "/v10.out"}, v10.mem);
        $writememh({DATA, "/v20.out"}, v20.mem);
        $writememh({DATA, "/w0.out"}, w0.mem);
        $writememh({DATA, "/x0.out"}, x0.mem);
        $writememh({DATA, "/y0.out"}, y0.mem);
        $writememh({DATA, "/z0.out"}, z0.mem);
    end
    logic [6:0] A0_0_addr0;
    logic [6:0] A0_0_addr1;
    logic [31:0] A0_0_write_data;
    logic A0_0_write_en;
    logic A0_0_clk;
    logic [31:0] A0_0_read_data;
    logic A0_0_done;
    logic [31:0] A_int_read0_0_in;
    logic A_int_read0_0_write_en;
    logic A_int_read0_0_clk;
    logic [31:0] A_int_read0_0_out;
    logic A_int_read0_0_done;
    logic [31:0] A_read0_0_in;
    logic A_read0_0_write_en;
    logic A_read0_0_clk;
    logic [31:0] A_read0_0_out;
    logic A_read0_0_done;
    logic [31:0] A_read1_0_in;
    logic A_read1_0_write_en;
    logic A_read1_0_clk;
    logic [31:0] A_read1_0_out;
    logic A_read1_0_done;
    logic [31:0] A_sh_read0_0_in;
    logic A_sh_read0_0_write_en;
    logic A_sh_read0_0_clk;
    logic [31:0] A_sh_read0_0_out;
    logic A_sh_read0_0_done;
    logic [6:0] add0_left;
    logic [6:0] add0_right;
    logic [6:0] add0_out;
    logic [6:0] add1_left;
    logic [6:0] add1_right;
    logic [6:0] add1_out;
    logic [31:0] add10_left;
    logic [31:0] add10_right;
    logic [31:0] add10_out;
    logic [31:0] alpha__0_in;
    logic alpha__0_write_en;
    logic alpha__0_clk;
    logic [31:0] alpha__0_out;
    logic alpha__0_done;
    logic [31:0] beta__0_in;
    logic beta__0_write_en;
    logic beta__0_clk;
    logic [31:0] beta__0_out;
    logic beta__0_done;
    logic [31:0] bin_read0_0_in;
    logic bin_read0_0_write_en;
    logic bin_read0_0_clk;
    logic [31:0] bin_read0_0_out;
    logic bin_read0_0_done;
    logic [31:0] bin_read1_0_in;
    logic bin_read1_0_write_en;
    logic bin_read1_0_clk;
    logic [31:0] bin_read1_0_out;
    logic bin_read1_0_done;
    logic [31:0] bin_read2_0_in;
    logic bin_read2_0_write_en;
    logic bin_read2_0_clk;
    logic [31:0] bin_read2_0_out;
    logic bin_read2_0_done;
    logic [31:0] bin_read3_0_in;
    logic bin_read3_0_write_en;
    logic bin_read3_0_clk;
    logic [31:0] bin_read3_0_out;
    logic bin_read3_0_done;
    logic [31:0] bin_read4_0_in;
    logic bin_read4_0_write_en;
    logic bin_read4_0_clk;
    logic [31:0] bin_read4_0_out;
    logic bin_read4_0_done;
    logic [31:0] bin_read5_0_in;
    logic bin_read5_0_write_en;
    logic bin_read5_0_clk;
    logic [31:0] bin_read5_0_out;
    logic bin_read5_0_done;
    logic const0_out;
    logic const1_out;
    logic [6:0] const10_out;
    logic [6:0] const11_out;
    logic [6:0] const12_out;
    logic [6:0] const13_out;
    logic [6:0] const14_out;
    logic [6:0] const16_out;
    logic [6:0] const19_out;
    logic [6:0] i0_in;
    logic i0_write_en;
    logic i0_clk;
    logic [6:0] i0_out;
    logic i0_done;
    logic [6:0] i1_in;
    logic i1_write_en;
    logic i1_clk;
    logic [6:0] i1_out;
    logic i1_done;
    logic [6:0] i2_in;
    logic i2_write_en;
    logic i2_clk;
    logic [6:0] i2_out;
    logic i2_done;
    logic [6:0] i3_in;
    logic i3_write_en;
    logic i3_clk;
    logic [6:0] i3_out;
    logic i3_done;
    logic [6:0] i4_in;
    logic i4_write_en;
    logic i4_clk;
    logic [6:0] i4_out;
    logic i4_done;
    logic [6:0] i5_in;
    logic i5_write_en;
    logic i5_clk;
    logic [6:0] i5_out;
    logic i5_done;
    logic [6:0] i6_in;
    logic i6_write_en;
    logic i6_clk;
    logic [6:0] i6_out;
    logic i6_done;
    logic [6:0] i7_in;
    logic i7_write_en;
    logic i7_clk;
    logic [6:0] i7_out;
    logic i7_done;
    logic [6:0] j0_in;
    logic j0_write_en;
    logic j0_clk;
    logic [6:0] j0_out;
    logic j0_done;
    logic [6:0] j1_in;
    logic j1_write_en;
    logic j1_clk;
    logic [6:0] j1_out;
    logic j1_done;
    logic [6:0] j2_in;
    logic j2_write_en;
    logic j2_clk;
    logic [6:0] j2_out;
    logic j2_done;
    logic [6:0] j3_in;
    logic j3_write_en;
    logic j3_clk;
    logic [6:0] j3_out;
    logic j3_done;
    logic [6:0] j4_in;
    logic j4_write_en;
    logic j4_clk;
    logic [6:0] j4_out;
    logic j4_done;
    logic [6:0] le0_left;
    logic [6:0] le0_right;
    logic le0_out;
    logic [6:0] le1_left;
    logic [6:0] le1_right;
    logic le1_out;
    logic [31:0] mult_pipe0_left;
    logic [31:0] mult_pipe0_right;
    logic mult_pipe0_go;
    logic mult_pipe0_clk;
    logic [31:0] mult_pipe0_out;
    logic mult_pipe0_done;
    logic [31:0] mult_pipe1_left;
    logic [31:0] mult_pipe1_right;
    logic mult_pipe1_go;
    logic mult_pipe1_clk;
    logic [31:0] mult_pipe1_out;
    logic mult_pipe1_done;
    logic [31:0] mult_pipe2_left;
    logic [31:0] mult_pipe2_right;
    logic mult_pipe2_go;
    logic mult_pipe2_clk;
    logic [31:0] mult_pipe2_out;
    logic mult_pipe2_done;
    logic [31:0] mult_pipe3_left;
    logic [31:0] mult_pipe3_right;
    logic mult_pipe3_go;
    logic mult_pipe3_clk;
    logic [31:0] mult_pipe3_out;
    logic mult_pipe3_done;
    logic [31:0] mult_pipe4_left;
    logic [31:0] mult_pipe4_right;
    logic mult_pipe4_go;
    logic mult_pipe4_clk;
    logic [31:0] mult_pipe4_out;
    logic mult_pipe4_done;
    logic [31:0] mult_pipe5_left;
    logic [31:0] mult_pipe5_right;
    logic mult_pipe5_go;
    logic mult_pipe5_clk;
    logic [31:0] mult_pipe5_out;
    logic mult_pipe5_done;
    logic [31:0] old_0_in;
    logic old_0_write_en;
    logic old_0_clk;
    logic [31:0] old_0_out;
    logic old_0_done;
    logic [31:0] old_1_in;
    logic old_1_write_en;
    logic old_1_clk;
    logic [31:0] old_1_out;
    logic old_1_done;
    logic [6:0] rsh0_left;
    logic [6:0] rsh0_right;
    logic [6:0] rsh0_out;
    logic [6:0] rsh1_left;
    logic [6:0] rsh1_right;
    logic [6:0] rsh1_out;
    logic [6:0] rsh10_left;
    logic [6:0] rsh10_right;
    logic [6:0] rsh10_out;
    logic [31:0] tmp1_0_in;
    logic tmp1_0_write_en;
    logic tmp1_0_clk;
    logic [31:0] tmp1_0_out;
    logic tmp1_0_done;
    logic [31:0] tmp2_0_in;
    logic tmp2_0_write_en;
    logic tmp2_0_clk;
    logic [31:0] tmp2_0_out;
    logic tmp2_0_done;
    logic [31:0] tmp3_0_in;
    logic tmp3_0_write_en;
    logic tmp3_0_clk;
    logic [31:0] tmp3_0_out;
    logic tmp3_0_done;
    logic [31:0] tmp4_0_in;
    logic tmp4_0_write_en;
    logic tmp4_0_clk;
    logic [31:0] tmp4_0_out;
    logic tmp4_0_done;
    logic [6:0] u10_addr0;
    logic [31:0] u10_write_data;
    logic u10_write_en;
    logic u10_clk;
    logic [31:0] u10_read_data;
    logic u10_done;
    logic [31:0] u1_int_read0_0_in;
    logic u1_int_read0_0_write_en;
    logic u1_int_read0_0_clk;
    logic [31:0] u1_int_read0_0_out;
    logic u1_int_read0_0_done;
    logic [31:0] u1_read0_0_in;
    logic u1_read0_0_write_en;
    logic u1_read0_0_clk;
    logic [31:0] u1_read0_0_out;
    logic u1_read0_0_done;
    logic [31:0] u1_sh_read0_0_in;
    logic u1_sh_read0_0_write_en;
    logic u1_sh_read0_0_clk;
    logic [31:0] u1_sh_read0_0_out;
    logic u1_sh_read0_0_done;
    logic [6:0] u20_addr0;
    logic [31:0] u20_write_data;
    logic u20_write_en;
    logic u20_clk;
    logic [31:0] u20_read_data;
    logic u20_done;
    logic [31:0] u2_int_read0_0_in;
    logic u2_int_read0_0_write_en;
    logic u2_int_read0_0_clk;
    logic [31:0] u2_int_read0_0_out;
    logic u2_int_read0_0_done;
    logic [31:0] u2_read0_0_in;
    logic u2_read0_0_write_en;
    logic u2_read0_0_clk;
    logic [31:0] u2_read0_0_out;
    logic u2_read0_0_done;
    logic [31:0] u2_sh_read0_0_in;
    logic u2_sh_read0_0_write_en;
    logic u2_sh_read0_0_clk;
    logic [31:0] u2_sh_read0_0_out;
    logic u2_sh_read0_0_done;
    logic [6:0] v10_addr0;
    logic [31:0] v10_write_data;
    logic v10_write_en;
    logic v10_clk;
    logic [31:0] v10_read_data;
    logic v10_done;
    logic [31:0] v1_int_read0_0_in;
    logic v1_int_read0_0_write_en;
    logic v1_int_read0_0_clk;
    logic [31:0] v1_int_read0_0_out;
    logic v1_int_read0_0_done;
    logic [31:0] v1_read0_0_in;
    logic v1_read0_0_write_en;
    logic v1_read0_0_clk;
    logic [31:0] v1_read0_0_out;
    logic v1_read0_0_done;
    logic [31:0] v1_sh_read0_0_in;
    logic v1_sh_read0_0_write_en;
    logic v1_sh_read0_0_clk;
    logic [31:0] v1_sh_read0_0_out;
    logic v1_sh_read0_0_done;
    logic [6:0] v20_addr0;
    logic [31:0] v20_write_data;
    logic v20_write_en;
    logic v20_clk;
    logic [31:0] v20_read_data;
    logic v20_done;
    logic [31:0] v2_int_read0_0_in;
    logic v2_int_read0_0_write_en;
    logic v2_int_read0_0_clk;
    logic [31:0] v2_int_read0_0_out;
    logic v2_int_read0_0_done;
    logic [31:0] v2_read0_0_in;
    logic v2_read0_0_write_en;
    logic v2_read0_0_clk;
    logic [31:0] v2_read0_0_out;
    logic v2_read0_0_done;
    logic [31:0] v2_sh_read0_0_in;
    logic v2_sh_read0_0_write_en;
    logic v2_sh_read0_0_clk;
    logic [31:0] v2_sh_read0_0_out;
    logic v2_sh_read0_0_done;
    logic [6:0] w0_addr0;
    logic [31:0] w0_write_data;
    logic w0_write_en;
    logic w0_clk;
    logic [31:0] w0_read_data;
    logic w0_done;
    logic [31:0] w_int_read0_0_in;
    logic w_int_read0_0_write_en;
    logic w_int_read0_0_clk;
    logic [31:0] w_int_read0_0_out;
    logic w_int_read0_0_done;
    logic [31:0] w_sh_read0_0_in;
    logic w_sh_read0_0_write_en;
    logic w_sh_read0_0_clk;
    logic [31:0] w_sh_read0_0_out;
    logic w_sh_read0_0_done;
    logic [6:0] x0_addr0;
    logic [31:0] x0_write_data;
    logic x0_write_en;
    logic x0_clk;
    logic [31:0] x0_read_data;
    logic x0_done;
    logic [31:0] x_int_read0_0_in;
    logic x_int_read0_0_write_en;
    logic x_int_read0_0_clk;
    logic [31:0] x_int_read0_0_out;
    logic x_int_read0_0_done;
    logic [31:0] x_read0_0_in;
    logic x_read0_0_write_en;
    logic x_read0_0_clk;
    logic [31:0] x_read0_0_out;
    logic x_read0_0_done;
    logic [31:0] x_sh_read0_0_in;
    logic x_sh_read0_0_write_en;
    logic x_sh_read0_0_clk;
    logic [31:0] x_sh_read0_0_out;
    logic x_sh_read0_0_done;
    logic [6:0] y0_addr0;
    logic [31:0] y0_write_data;
    logic y0_write_en;
    logic y0_clk;
    logic [31:0] y0_read_data;
    logic y0_done;
    logic [31:0] y_int_read0_0_in;
    logic y_int_read0_0_write_en;
    logic y_int_read0_0_clk;
    logic [31:0] y_int_read0_0_out;
    logic y_int_read0_0_done;
    logic [31:0] y_read0_0_in;
    logic y_read0_0_write_en;
    logic y_read0_0_clk;
    logic [31:0] y_read0_0_out;
    logic y_read0_0_done;
    logic [31:0] y_sh_read0_0_in;
    logic y_sh_read0_0_write_en;
    logic y_sh_read0_0_clk;
    logic [31:0] y_sh_read0_0_out;
    logic y_sh_read0_0_done;
    logic [6:0] z0_addr0;
    logic [31:0] z0_write_data;
    logic z0_write_en;
    logic z0_clk;
    logic [31:0] z0_read_data;
    logic z0_done;
    logic [31:0] z_int_read0_0_in;
    logic z_int_read0_0_write_en;
    logic z_int_read0_0_clk;
    logic [31:0] z_int_read0_0_out;
    logic z_int_read0_0_done;
    logic [31:0] z_sh_read0_0_in;
    logic z_sh_read0_0_write_en;
    logic z_sh_read0_0_clk;
    logic [31:0] z_sh_read0_0_out;
    logic z_sh_read0_0_done;
    logic par_reset_in;
    logic par_reset_write_en;
    logic par_reset_clk;
    logic par_reset_out;
    logic par_reset_done;
    logic par_done_reg_in;
    logic par_done_reg_write_en;
    logic par_done_reg_clk;
    logic par_done_reg_out;
    logic par_done_reg_done;
    logic par_done_reg0_in;
    logic par_done_reg0_write_en;
    logic par_done_reg0_clk;
    logic par_done_reg0_out;
    logic par_done_reg0_done;
    logic par_reset0_in;
    logic par_reset0_write_en;
    logic par_reset0_clk;
    logic par_reset0_out;
    logic par_reset0_done;
    logic par_done_reg1_in;
    logic par_done_reg1_write_en;
    logic par_done_reg1_clk;
    logic par_done_reg1_out;
    logic par_done_reg1_done;
    logic par_done_reg2_in;
    logic par_done_reg2_write_en;
    logic par_done_reg2_clk;
    logic par_done_reg2_out;
    logic par_done_reg2_done;
    logic par_reset1_in;
    logic par_reset1_write_en;
    logic par_reset1_clk;
    logic par_reset1_out;
    logic par_reset1_done;
    logic par_done_reg3_in;
    logic par_done_reg3_write_en;
    logic par_done_reg3_clk;
    logic par_done_reg3_out;
    logic par_done_reg3_done;
    logic par_done_reg4_in;
    logic par_done_reg4_write_en;
    logic par_done_reg4_clk;
    logic par_done_reg4_out;
    logic par_done_reg4_done;
    logic par_reset2_in;
    logic par_reset2_write_en;
    logic par_reset2_clk;
    logic par_reset2_out;
    logic par_reset2_done;
    logic par_done_reg5_in;
    logic par_done_reg5_write_en;
    logic par_done_reg5_clk;
    logic par_done_reg5_out;
    logic par_done_reg5_done;
    logic par_done_reg6_in;
    logic par_done_reg6_write_en;
    logic par_done_reg6_clk;
    logic par_done_reg6_out;
    logic par_done_reg6_done;
    logic par_reset3_in;
    logic par_reset3_write_en;
    logic par_reset3_clk;
    logic par_reset3_out;
    logic par_reset3_done;
    logic par_done_reg7_in;
    logic par_done_reg7_write_en;
    logic par_done_reg7_clk;
    logic par_done_reg7_out;
    logic par_done_reg7_done;
    logic par_done_reg8_in;
    logic par_done_reg8_write_en;
    logic par_done_reg8_clk;
    logic par_done_reg8_out;
    logic par_done_reg8_done;
    logic par_reset4_in;
    logic par_reset4_write_en;
    logic par_reset4_clk;
    logic par_reset4_out;
    logic par_reset4_done;
    logic par_done_reg9_in;
    logic par_done_reg9_write_en;
    logic par_done_reg9_clk;
    logic par_done_reg9_out;
    logic par_done_reg9_done;
    logic par_done_reg10_in;
    logic par_done_reg10_write_en;
    logic par_done_reg10_clk;
    logic par_done_reg10_out;
    logic par_done_reg10_done;
    logic par_reset5_in;
    logic par_reset5_write_en;
    logic par_reset5_clk;
    logic par_reset5_out;
    logic par_reset5_done;
    logic par_done_reg11_in;
    logic par_done_reg11_write_en;
    logic par_done_reg11_clk;
    logic par_done_reg11_out;
    logic par_done_reg11_done;
    logic par_done_reg12_in;
    logic par_done_reg12_write_en;
    logic par_done_reg12_clk;
    logic par_done_reg12_out;
    logic par_done_reg12_done;
    logic [31:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic [31:0] fsm_out;
    logic fsm_done;
    logic cond_computed_in;
    logic cond_computed_write_en;
    logic cond_computed_clk;
    logic cond_computed_out;
    logic cond_computed_done;
    logic cond_stored_in;
    logic cond_stored_write_en;
    logic cond_stored_clk;
    logic cond_stored_out;
    logic cond_stored_done;
    logic done_reg_in;
    logic done_reg_write_en;
    logic done_reg_clk;
    logic done_reg_out;
    logic done_reg_done;
    logic [31:0] fsm0_in;
    logic fsm0_write_en;
    logic fsm0_clk;
    logic [31:0] fsm0_out;
    logic fsm0_done;
    logic [31:0] fsm1_in;
    logic fsm1_write_en;
    logic fsm1_clk;
    logic [31:0] fsm1_out;
    logic fsm1_done;
    logic cond_computed0_in;
    logic cond_computed0_write_en;
    logic cond_computed0_clk;
    logic cond_computed0_out;
    logic cond_computed0_done;
    logic cond_stored0_in;
    logic cond_stored0_write_en;
    logic cond_stored0_clk;
    logic cond_stored0_out;
    logic cond_stored0_done;
    logic done_reg0_in;
    logic done_reg0_write_en;
    logic done_reg0_clk;
    logic done_reg0_out;
    logic done_reg0_done;
    logic [31:0] fsm2_in;
    logic fsm2_write_en;
    logic fsm2_clk;
    logic [31:0] fsm2_out;
    logic fsm2_done;
    logic cond_computed1_in;
    logic cond_computed1_write_en;
    logic cond_computed1_clk;
    logic cond_computed1_out;
    logic cond_computed1_done;
    logic cond_stored1_in;
    logic cond_stored1_write_en;
    logic cond_stored1_clk;
    logic cond_stored1_out;
    logic cond_stored1_done;
    logic done_reg1_in;
    logic done_reg1_write_en;
    logic done_reg1_clk;
    logic done_reg1_out;
    logic done_reg1_done;
    logic [31:0] fsm3_in;
    logic fsm3_write_en;
    logic fsm3_clk;
    logic [31:0] fsm3_out;
    logic fsm3_done;
    logic par_reset6_in;
    logic par_reset6_write_en;
    logic par_reset6_clk;
    logic par_reset6_out;
    logic par_reset6_done;
    logic par_done_reg13_in;
    logic par_done_reg13_write_en;
    logic par_done_reg13_clk;
    logic par_done_reg13_out;
    logic par_done_reg13_done;
    logic par_done_reg14_in;
    logic par_done_reg14_write_en;
    logic par_done_reg14_clk;
    logic par_done_reg14_out;
    logic par_done_reg14_done;
    logic par_done_reg15_in;
    logic par_done_reg15_write_en;
    logic par_done_reg15_clk;
    logic par_done_reg15_out;
    logic par_done_reg15_done;
    logic par_done_reg16_in;
    logic par_done_reg16_write_en;
    logic par_done_reg16_clk;
    logic par_done_reg16_out;
    logic par_done_reg16_done;
    logic par_reset7_in;
    logic par_reset7_write_en;
    logic par_reset7_clk;
    logic par_reset7_out;
    logic par_reset7_done;
    logic par_done_reg17_in;
    logic par_done_reg17_write_en;
    logic par_done_reg17_clk;
    logic par_done_reg17_out;
    logic par_done_reg17_done;
    logic par_done_reg18_in;
    logic par_done_reg18_write_en;
    logic par_done_reg18_clk;
    logic par_done_reg18_out;
    logic par_done_reg18_done;
    logic par_done_reg19_in;
    logic par_done_reg19_write_en;
    logic par_done_reg19_clk;
    logic par_done_reg19_out;
    logic par_done_reg19_done;
    logic par_done_reg20_in;
    logic par_done_reg20_write_en;
    logic par_done_reg20_clk;
    logic par_done_reg20_out;
    logic par_done_reg20_done;
    logic [31:0] fsm4_in;
    logic fsm4_write_en;
    logic fsm4_clk;
    logic [31:0] fsm4_out;
    logic fsm4_done;
    logic par_reset8_in;
    logic par_reset8_write_en;
    logic par_reset8_clk;
    logic par_reset8_out;
    logic par_reset8_done;
    logic par_done_reg21_in;
    logic par_done_reg21_write_en;
    logic par_done_reg21_clk;
    logic par_done_reg21_out;
    logic par_done_reg21_done;
    logic par_done_reg22_in;
    logic par_done_reg22_write_en;
    logic par_done_reg22_clk;
    logic par_done_reg22_out;
    logic par_done_reg22_done;
    logic [31:0] fsm5_in;
    logic fsm5_write_en;
    logic fsm5_clk;
    logic [31:0] fsm5_out;
    logic fsm5_done;
    logic cond_computed2_in;
    logic cond_computed2_write_en;
    logic cond_computed2_clk;
    logic cond_computed2_out;
    logic cond_computed2_done;
    logic cond_stored2_in;
    logic cond_stored2_write_en;
    logic cond_stored2_clk;
    logic cond_stored2_out;
    logic cond_stored2_done;
    logic done_reg2_in;
    logic done_reg2_write_en;
    logic done_reg2_clk;
    logic done_reg2_out;
    logic done_reg2_done;
    logic [31:0] fsm6_in;
    logic fsm6_write_en;
    logic fsm6_clk;
    logic [31:0] fsm6_out;
    logic fsm6_done;
    logic cond_computed3_in;
    logic cond_computed3_write_en;
    logic cond_computed3_clk;
    logic cond_computed3_out;
    logic cond_computed3_done;
    logic cond_stored3_in;
    logic cond_stored3_write_en;
    logic cond_stored3_clk;
    logic cond_stored3_out;
    logic cond_stored3_done;
    logic done_reg3_in;
    logic done_reg3_write_en;
    logic done_reg3_clk;
    logic done_reg3_out;
    logic done_reg3_done;
    logic par_reset9_in;
    logic par_reset9_write_en;
    logic par_reset9_clk;
    logic par_reset9_out;
    logic par_reset9_done;
    logic par_done_reg23_in;
    logic par_done_reg23_write_en;
    logic par_done_reg23_clk;
    logic par_done_reg23_out;
    logic par_done_reg23_done;
    logic par_done_reg24_in;
    logic par_done_reg24_write_en;
    logic par_done_reg24_clk;
    logic par_done_reg24_out;
    logic par_done_reg24_done;
    logic [31:0] fsm7_in;
    logic fsm7_write_en;
    logic fsm7_clk;
    logic [31:0] fsm7_out;
    logic fsm7_done;
    logic cond_computed4_in;
    logic cond_computed4_write_en;
    logic cond_computed4_clk;
    logic cond_computed4_out;
    logic cond_computed4_done;
    logic cond_stored4_in;
    logic cond_stored4_write_en;
    logic cond_stored4_clk;
    logic cond_stored4_out;
    logic cond_stored4_done;
    logic done_reg4_in;
    logic done_reg4_write_en;
    logic done_reg4_clk;
    logic done_reg4_out;
    logic done_reg4_done;
    logic [31:0] fsm8_in;
    logic fsm8_write_en;
    logic fsm8_clk;
    logic [31:0] fsm8_out;
    logic fsm8_done;
    logic cond_computed5_in;
    logic cond_computed5_write_en;
    logic cond_computed5_clk;
    logic cond_computed5_out;
    logic cond_computed5_done;
    logic cond_stored5_in;
    logic cond_stored5_write_en;
    logic cond_stored5_clk;
    logic cond_stored5_out;
    logic cond_stored5_done;
    logic done_reg5_in;
    logic done_reg5_write_en;
    logic done_reg5_clk;
    logic done_reg5_out;
    logic done_reg5_done;
    logic par_reset10_in;
    logic par_reset10_write_en;
    logic par_reset10_clk;
    logic par_reset10_out;
    logic par_reset10_done;
    logic par_done_reg25_in;
    logic par_done_reg25_write_en;
    logic par_done_reg25_clk;
    logic par_done_reg25_out;
    logic par_done_reg25_done;
    logic par_done_reg26_in;
    logic par_done_reg26_write_en;
    logic par_done_reg26_clk;
    logic par_done_reg26_out;
    logic par_done_reg26_done;
    logic [31:0] fsm9_in;
    logic fsm9_write_en;
    logic fsm9_clk;
    logic [31:0] fsm9_out;
    logic fsm9_done;
    logic cond_computed6_in;
    logic cond_computed6_write_en;
    logic cond_computed6_clk;
    logic cond_computed6_out;
    logic cond_computed6_done;
    logic cond_stored6_in;
    logic cond_stored6_write_en;
    logic cond_stored6_clk;
    logic cond_stored6_out;
    logic cond_stored6_done;
    logic done_reg6_in;
    logic done_reg6_write_en;
    logic done_reg6_clk;
    logic done_reg6_out;
    logic done_reg6_done;
    logic par_reset11_in;
    logic par_reset11_write_en;
    logic par_reset11_clk;
    logic par_reset11_out;
    logic par_reset11_done;
    logic par_done_reg27_in;
    logic par_done_reg27_write_en;
    logic par_done_reg27_clk;
    logic par_done_reg27_out;
    logic par_done_reg27_done;
    logic par_done_reg28_in;
    logic par_done_reg28_write_en;
    logic par_done_reg28_clk;
    logic par_done_reg28_out;
    logic par_done_reg28_done;
    logic [31:0] fsm10_in;
    logic fsm10_write_en;
    logic fsm10_clk;
    logic [31:0] fsm10_out;
    logic fsm10_done;
    logic cond_computed7_in;
    logic cond_computed7_write_en;
    logic cond_computed7_clk;
    logic cond_computed7_out;
    logic cond_computed7_done;
    logic cond_stored7_in;
    logic cond_stored7_write_en;
    logic cond_stored7_clk;
    logic cond_stored7_out;
    logic cond_stored7_done;
    logic done_reg7_in;
    logic done_reg7_write_en;
    logic done_reg7_clk;
    logic done_reg7_out;
    logic done_reg7_done;
    logic [31:0] fsm11_in;
    logic fsm11_write_en;
    logic fsm11_clk;
    logic [31:0] fsm11_out;
    logic fsm11_done;
    logic cond_computed8_in;
    logic cond_computed8_write_en;
    logic cond_computed8_clk;
    logic cond_computed8_out;
    logic cond_computed8_done;
    logic cond_stored8_in;
    logic cond_stored8_write_en;
    logic cond_stored8_clk;
    logic cond_stored8_out;
    logic cond_stored8_done;
    logic done_reg8_in;
    logic done_reg8_write_en;
    logic done_reg8_clk;
    logic done_reg8_out;
    logic done_reg8_done;
    logic par_reset12_in;
    logic par_reset12_write_en;
    logic par_reset12_clk;
    logic par_reset12_out;
    logic par_reset12_done;
    logic par_done_reg29_in;
    logic par_done_reg29_write_en;
    logic par_done_reg29_clk;
    logic par_done_reg29_out;
    logic par_done_reg29_done;
    logic par_done_reg30_in;
    logic par_done_reg30_write_en;
    logic par_done_reg30_clk;
    logic par_done_reg30_out;
    logic par_done_reg30_done;
    logic par_reset13_in;
    logic par_reset13_write_en;
    logic par_reset13_clk;
    logic par_reset13_out;
    logic par_reset13_done;
    logic par_done_reg31_in;
    logic par_done_reg31_write_en;
    logic par_done_reg31_clk;
    logic par_done_reg31_out;
    logic par_done_reg31_done;
    logic par_done_reg32_in;
    logic par_done_reg32_write_en;
    logic par_done_reg32_clk;
    logic par_done_reg32_out;
    logic par_done_reg32_done;
    logic par_reset14_in;
    logic par_reset14_write_en;
    logic par_reset14_clk;
    logic par_reset14_out;
    logic par_reset14_done;
    logic par_done_reg33_in;
    logic par_done_reg33_write_en;
    logic par_done_reg33_clk;
    logic par_done_reg33_out;
    logic par_done_reg33_done;
    logic par_done_reg34_in;
    logic par_done_reg34_write_en;
    logic par_done_reg34_clk;
    logic par_done_reg34_out;
    logic par_done_reg34_done;
    logic par_reset15_in;
    logic par_reset15_write_en;
    logic par_reset15_clk;
    logic par_reset15_out;
    logic par_reset15_done;
    logic par_done_reg35_in;
    logic par_done_reg35_write_en;
    logic par_done_reg35_clk;
    logic par_done_reg35_out;
    logic par_done_reg35_done;
    logic par_done_reg36_in;
    logic par_done_reg36_write_en;
    logic par_done_reg36_clk;
    logic par_done_reg36_out;
    logic par_done_reg36_done;
    logic par_reset16_in;
    logic par_reset16_write_en;
    logic par_reset16_clk;
    logic par_reset16_out;
    logic par_reset16_done;
    logic par_done_reg37_in;
    logic par_done_reg37_write_en;
    logic par_done_reg37_clk;
    logic par_done_reg37_out;
    logic par_done_reg37_done;
    logic par_done_reg38_in;
    logic par_done_reg38_write_en;
    logic par_done_reg38_clk;
    logic par_done_reg38_out;
    logic par_done_reg38_done;
    logic par_reset17_in;
    logic par_reset17_write_en;
    logic par_reset17_clk;
    logic par_reset17_out;
    logic par_reset17_done;
    logic par_done_reg39_in;
    logic par_done_reg39_write_en;
    logic par_done_reg39_clk;
    logic par_done_reg39_out;
    logic par_done_reg39_done;
    logic par_done_reg40_in;
    logic par_done_reg40_write_en;
    logic par_done_reg40_clk;
    logic par_done_reg40_out;
    logic par_done_reg40_done;
    logic par_reset18_in;
    logic par_reset18_write_en;
    logic par_reset18_clk;
    logic par_reset18_out;
    logic par_reset18_done;
    logic par_done_reg41_in;
    logic par_done_reg41_write_en;
    logic par_done_reg41_clk;
    logic par_done_reg41_out;
    logic par_done_reg41_done;
    logic par_done_reg42_in;
    logic par_done_reg42_write_en;
    logic par_done_reg42_clk;
    logic par_done_reg42_out;
    logic par_done_reg42_done;
    logic [31:0] fsm12_in;
    logic fsm12_write_en;
    logic fsm12_clk;
    logic [31:0] fsm12_out;
    logic fsm12_done;
    logic cond_computed9_in;
    logic cond_computed9_write_en;
    logic cond_computed9_clk;
    logic cond_computed9_out;
    logic cond_computed9_done;
    logic cond_stored9_in;
    logic cond_stored9_write_en;
    logic cond_stored9_clk;
    logic cond_stored9_out;
    logic cond_stored9_done;
    logic done_reg9_in;
    logic done_reg9_write_en;
    logic done_reg9_clk;
    logic done_reg9_out;
    logic done_reg9_done;
    logic [31:0] fsm13_in;
    logic fsm13_write_en;
    logic fsm13_clk;
    logic [31:0] fsm13_out;
    logic fsm13_done;
    logic [31:0] fsm14_in;
    logic fsm14_write_en;
    logic fsm14_clk;
    logic [31:0] fsm14_out;
    logic fsm14_done;
    logic cond_computed10_in;
    logic cond_computed10_write_en;
    logic cond_computed10_clk;
    logic cond_computed10_out;
    logic cond_computed10_done;
    logic cond_stored10_in;
    logic cond_stored10_write_en;
    logic cond_stored10_clk;
    logic cond_stored10_out;
    logic cond_stored10_done;
    logic done_reg10_in;
    logic done_reg10_write_en;
    logic done_reg10_clk;
    logic done_reg10_out;
    logic done_reg10_done;
    logic [31:0] fsm15_in;
    logic fsm15_write_en;
    logic fsm15_clk;
    logic [31:0] fsm15_out;
    logic fsm15_done;
    logic cond_computed11_in;
    logic cond_computed11_write_en;
    logic cond_computed11_clk;
    logic cond_computed11_out;
    logic cond_computed11_done;
    logic cond_stored11_in;
    logic cond_stored11_write_en;
    logic cond_stored11_clk;
    logic cond_stored11_out;
    logic cond_stored11_done;
    logic done_reg11_in;
    logic done_reg11_write_en;
    logic done_reg11_clk;
    logic done_reg11_out;
    logic done_reg11_done;
    logic [31:0] fsm16_in;
    logic fsm16_write_en;
    logic fsm16_clk;
    logic [31:0] fsm16_out;
    logic fsm16_done;
    logic par_reset19_in;
    logic par_reset19_write_en;
    logic par_reset19_clk;
    logic par_reset19_out;
    logic par_reset19_done;
    logic par_done_reg43_in;
    logic par_done_reg43_write_en;
    logic par_done_reg43_clk;
    logic par_done_reg43_out;
    logic par_done_reg43_done;
    logic par_done_reg44_in;
    logic par_done_reg44_write_en;
    logic par_done_reg44_clk;
    logic par_done_reg44_out;
    logic par_done_reg44_done;
    logic [31:0] fsm17_in;
    logic fsm17_write_en;
    logic fsm17_clk;
    logic [31:0] fsm17_out;
    logic fsm17_done;
    std_mem_d2 # (
        .d0_idx_size(7),
        .d0_size(64),
        .d1_idx_size(7),
        .d1_size(64),
        .width(32)
    ) A0_0 (
        .addr0(A0_0_addr0),
        .addr1(A0_0_addr1),
        .clk(A0_0_clk),
        .done(A0_0_done),
        .read_data(A0_0_read_data),
        .write_data(A0_0_write_data),
        .write_en(A0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_int_read0_0 (
        .clk(A_int_read0_0_clk),
        .done(A_int_read0_0_done),
        .in(A_int_read0_0_in),
        .out(A_int_read0_0_out),
        .write_en(A_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_read0_0 (
        .clk(A_read0_0_clk),
        .done(A_read0_0_done),
        .in(A_read0_0_in),
        .out(A_read0_0_out),
        .write_en(A_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_read1_0 (
        .clk(A_read1_0_clk),
        .done(A_read1_0_done),
        .in(A_read1_0_in),
        .out(A_read1_0_out),
        .write_en(A_read1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_sh_read0_0 (
        .clk(A_sh_read0_0_clk),
        .done(A_sh_read0_0_done),
        .in(A_sh_read0_0_in),
        .out(A_sh_read0_0_out),
        .write_en(A_sh_read0_0_write_en)
    );
    std_add # (
        .width(7)
    ) add0 (
        .left(add0_left),
        .out(add0_out),
        .right(add0_right)
    );
    std_add # (
        .width(7)
    ) add1 (
        .left(add1_left),
        .out(add1_out),
        .right(add1_right)
    );
    std_add # (
        .width(32)
    ) add10 (
        .left(add10_left),
        .out(add10_out),
        .right(add10_right)
    );
    std_reg # (
        .width(32)
    ) alpha__0 (
        .clk(alpha__0_clk),
        .done(alpha__0_done),
        .in(alpha__0_in),
        .out(alpha__0_out),
        .write_en(alpha__0_write_en)
    );
    std_reg # (
        .width(32)
    ) beta__0 (
        .clk(beta__0_clk),
        .done(beta__0_done),
        .in(beta__0_in),
        .out(beta__0_out),
        .write_en(beta__0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read0_0 (
        .clk(bin_read0_0_clk),
        .done(bin_read0_0_done),
        .in(bin_read0_0_in),
        .out(bin_read0_0_out),
        .write_en(bin_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read1_0 (
        .clk(bin_read1_0_clk),
        .done(bin_read1_0_done),
        .in(bin_read1_0_in),
        .out(bin_read1_0_out),
        .write_en(bin_read1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read2_0 (
        .clk(bin_read2_0_clk),
        .done(bin_read2_0_done),
        .in(bin_read2_0_in),
        .out(bin_read2_0_out),
        .write_en(bin_read2_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read3_0 (
        .clk(bin_read3_0_clk),
        .done(bin_read3_0_done),
        .in(bin_read3_0_in),
        .out(bin_read3_0_out),
        .write_en(bin_read3_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read4_0 (
        .clk(bin_read4_0_clk),
        .done(bin_read4_0_done),
        .in(bin_read4_0_in),
        .out(bin_read4_0_out),
        .write_en(bin_read4_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read5_0 (
        .clk(bin_read5_0_clk),
        .done(bin_read5_0_done),
        .in(bin_read5_0_in),
        .out(bin_read5_0_out),
        .write_en(bin_read5_0_write_en)
    );
    std_const # (
        .value(0),
        .width(1)
    ) const0 (
        .out(const0_out)
    );
    std_const # (
        .value(0),
        .width(1)
    ) const1 (
        .out(const1_out)
    );
    std_const # (
        .value(0),
        .width(7)
    ) const10 (
        .out(const10_out)
    );
    std_const # (
        .value(0),
        .width(7)
    ) const11 (
        .out(const11_out)
    );
    std_const # (
        .value(1),
        .width(7)
    ) const12 (
        .out(const12_out)
    );
    std_const # (
        .value(0),
        .width(7)
    ) const13 (
        .out(const13_out)
    );
    std_const # (
        .value(63),
        .width(7)
    ) const14 (
        .out(const14_out)
    );
    std_const # (
        .value(63),
        .width(7)
    ) const16 (
        .out(const16_out)
    );
    std_const # (
        .value(1),
        .width(7)
    ) const19 (
        .out(const19_out)
    );
    std_reg # (
        .width(7)
    ) i0 (
        .clk(i0_clk),
        .done(i0_done),
        .in(i0_in),
        .out(i0_out),
        .write_en(i0_write_en)
    );
    std_reg # (
        .width(7)
    ) i1 (
        .clk(i1_clk),
        .done(i1_done),
        .in(i1_in),
        .out(i1_out),
        .write_en(i1_write_en)
    );
    std_reg # (
        .width(7)
    ) i2 (
        .clk(i2_clk),
        .done(i2_done),
        .in(i2_in),
        .out(i2_out),
        .write_en(i2_write_en)
    );
    std_reg # (
        .width(7)
    ) i3 (
        .clk(i3_clk),
        .done(i3_done),
        .in(i3_in),
        .out(i3_out),
        .write_en(i3_write_en)
    );
    std_reg # (
        .width(7)
    ) i4 (
        .clk(i4_clk),
        .done(i4_done),
        .in(i4_in),
        .out(i4_out),
        .write_en(i4_write_en)
    );
    std_reg # (
        .width(7)
    ) i5 (
        .clk(i5_clk),
        .done(i5_done),
        .in(i5_in),
        .out(i5_out),
        .write_en(i5_write_en)
    );
    std_reg # (
        .width(7)
    ) i6 (
        .clk(i6_clk),
        .done(i6_done),
        .in(i6_in),
        .out(i6_out),
        .write_en(i6_write_en)
    );
    std_reg # (
        .width(7)
    ) i7 (
        .clk(i7_clk),
        .done(i7_done),
        .in(i7_in),
        .out(i7_out),
        .write_en(i7_write_en)
    );
    std_reg # (
        .width(7)
    ) j0 (
        .clk(j0_clk),
        .done(j0_done),
        .in(j0_in),
        .out(j0_out),
        .write_en(j0_write_en)
    );
    std_reg # (
        .width(7)
    ) j1 (
        .clk(j1_clk),
        .done(j1_done),
        .in(j1_in),
        .out(j1_out),
        .write_en(j1_write_en)
    );
    std_reg # (
        .width(7)
    ) j2 (
        .clk(j2_clk),
        .done(j2_done),
        .in(j2_in),
        .out(j2_out),
        .write_en(j2_write_en)
    );
    std_reg # (
        .width(7)
    ) j3 (
        .clk(j3_clk),
        .done(j3_done),
        .in(j3_in),
        .out(j3_out),
        .write_en(j3_write_en)
    );
    std_reg # (
        .width(7)
    ) j4 (
        .clk(j4_clk),
        .done(j4_done),
        .in(j4_in),
        .out(j4_out),
        .write_en(j4_write_en)
    );
    std_le # (
        .width(7)
    ) le0 (
        .left(le0_left),
        .out(le0_out),
        .right(le0_right)
    );
    std_le # (
        .width(7)
    ) le1 (
        .left(le1_left),
        .out(le1_out),
        .right(le1_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe0 (
        .clk(mult_pipe0_clk),
        .done(mult_pipe0_done),
        .go(mult_pipe0_go),
        .left(mult_pipe0_left),
        .out(mult_pipe0_out),
        .right(mult_pipe0_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe1 (
        .clk(mult_pipe1_clk),
        .done(mult_pipe1_done),
        .go(mult_pipe1_go),
        .left(mult_pipe1_left),
        .out(mult_pipe1_out),
        .right(mult_pipe1_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe2 (
        .clk(mult_pipe2_clk),
        .done(mult_pipe2_done),
        .go(mult_pipe2_go),
        .left(mult_pipe2_left),
        .out(mult_pipe2_out),
        .right(mult_pipe2_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe3 (
        .clk(mult_pipe3_clk),
        .done(mult_pipe3_done),
        .go(mult_pipe3_go),
        .left(mult_pipe3_left),
        .out(mult_pipe3_out),
        .right(mult_pipe3_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe4 (
        .clk(mult_pipe4_clk),
        .done(mult_pipe4_done),
        .go(mult_pipe4_go),
        .left(mult_pipe4_left),
        .out(mult_pipe4_out),
        .right(mult_pipe4_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe5 (
        .clk(mult_pipe5_clk),
        .done(mult_pipe5_done),
        .go(mult_pipe5_go),
        .left(mult_pipe5_left),
        .out(mult_pipe5_out),
        .right(mult_pipe5_right)
    );
    std_reg # (
        .width(32)
    ) old_0 (
        .clk(old_0_clk),
        .done(old_0_done),
        .in(old_0_in),
        .out(old_0_out),
        .write_en(old_0_write_en)
    );
    std_reg # (
        .width(32)
    ) old_1 (
        .clk(old_1_clk),
        .done(old_1_done),
        .in(old_1_in),
        .out(old_1_out),
        .write_en(old_1_write_en)
    );
    std_rsh # (
        .width(7)
    ) rsh0 (
        .left(rsh0_left),
        .out(rsh0_out),
        .right(rsh0_right)
    );
    std_rsh # (
        .width(7)
    ) rsh1 (
        .left(rsh1_left),
        .out(rsh1_out),
        .right(rsh1_right)
    );
    std_rsh # (
        .width(7)
    ) rsh10 (
        .left(rsh10_left),
        .out(rsh10_out),
        .right(rsh10_right)
    );
    std_reg # (
        .width(32)
    ) tmp1_0 (
        .clk(tmp1_0_clk),
        .done(tmp1_0_done),
        .in(tmp1_0_in),
        .out(tmp1_0_out),
        .write_en(tmp1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) tmp2_0 (
        .clk(tmp2_0_clk),
        .done(tmp2_0_done),
        .in(tmp2_0_in),
        .out(tmp2_0_out),
        .write_en(tmp2_0_write_en)
    );
    std_reg # (
        .width(32)
    ) tmp3_0 (
        .clk(tmp3_0_clk),
        .done(tmp3_0_done),
        .in(tmp3_0_in),
        .out(tmp3_0_out),
        .write_en(tmp3_0_write_en)
    );
    std_reg # (
        .width(32)
    ) tmp4_0 (
        .clk(tmp4_0_clk),
        .done(tmp4_0_done),
        .in(tmp4_0_in),
        .out(tmp4_0_out),
        .write_en(tmp4_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) u10 (
        .addr0(u10_addr0),
        .clk(u10_clk),
        .done(u10_done),
        .read_data(u10_read_data),
        .write_data(u10_write_data),
        .write_en(u10_write_en)
    );
    std_reg # (
        .width(32)
    ) u1_int_read0_0 (
        .clk(u1_int_read0_0_clk),
        .done(u1_int_read0_0_done),
        .in(u1_int_read0_0_in),
        .out(u1_int_read0_0_out),
        .write_en(u1_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) u1_read0_0 (
        .clk(u1_read0_0_clk),
        .done(u1_read0_0_done),
        .in(u1_read0_0_in),
        .out(u1_read0_0_out),
        .write_en(u1_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) u1_sh_read0_0 (
        .clk(u1_sh_read0_0_clk),
        .done(u1_sh_read0_0_done),
        .in(u1_sh_read0_0_in),
        .out(u1_sh_read0_0_out),
        .write_en(u1_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) u20 (
        .addr0(u20_addr0),
        .clk(u20_clk),
        .done(u20_done),
        .read_data(u20_read_data),
        .write_data(u20_write_data),
        .write_en(u20_write_en)
    );
    std_reg # (
        .width(32)
    ) u2_int_read0_0 (
        .clk(u2_int_read0_0_clk),
        .done(u2_int_read0_0_done),
        .in(u2_int_read0_0_in),
        .out(u2_int_read0_0_out),
        .write_en(u2_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) u2_read0_0 (
        .clk(u2_read0_0_clk),
        .done(u2_read0_0_done),
        .in(u2_read0_0_in),
        .out(u2_read0_0_out),
        .write_en(u2_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) u2_sh_read0_0 (
        .clk(u2_sh_read0_0_clk),
        .done(u2_sh_read0_0_done),
        .in(u2_sh_read0_0_in),
        .out(u2_sh_read0_0_out),
        .write_en(u2_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) v10 (
        .addr0(v10_addr0),
        .clk(v10_clk),
        .done(v10_done),
        .read_data(v10_read_data),
        .write_data(v10_write_data),
        .write_en(v10_write_en)
    );
    std_reg # (
        .width(32)
    ) v1_int_read0_0 (
        .clk(v1_int_read0_0_clk),
        .done(v1_int_read0_0_done),
        .in(v1_int_read0_0_in),
        .out(v1_int_read0_0_out),
        .write_en(v1_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) v1_read0_0 (
        .clk(v1_read0_0_clk),
        .done(v1_read0_0_done),
        .in(v1_read0_0_in),
        .out(v1_read0_0_out),
        .write_en(v1_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) v1_sh_read0_0 (
        .clk(v1_sh_read0_0_clk),
        .done(v1_sh_read0_0_done),
        .in(v1_sh_read0_0_in),
        .out(v1_sh_read0_0_out),
        .write_en(v1_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) v20 (
        .addr0(v20_addr0),
        .clk(v20_clk),
        .done(v20_done),
        .read_data(v20_read_data),
        .write_data(v20_write_data),
        .write_en(v20_write_en)
    );
    std_reg # (
        .width(32)
    ) v2_int_read0_0 (
        .clk(v2_int_read0_0_clk),
        .done(v2_int_read0_0_done),
        .in(v2_int_read0_0_in),
        .out(v2_int_read0_0_out),
        .write_en(v2_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) v2_read0_0 (
        .clk(v2_read0_0_clk),
        .done(v2_read0_0_done),
        .in(v2_read0_0_in),
        .out(v2_read0_0_out),
        .write_en(v2_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) v2_sh_read0_0 (
        .clk(v2_sh_read0_0_clk),
        .done(v2_sh_read0_0_done),
        .in(v2_sh_read0_0_in),
        .out(v2_sh_read0_0_out),
        .write_en(v2_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) w0 (
        .addr0(w0_addr0),
        .clk(w0_clk),
        .done(w0_done),
        .read_data(w0_read_data),
        .write_data(w0_write_data),
        .write_en(w0_write_en)
    );
    std_reg # (
        .width(32)
    ) w_int_read0_0 (
        .clk(w_int_read0_0_clk),
        .done(w_int_read0_0_done),
        .in(w_int_read0_0_in),
        .out(w_int_read0_0_out),
        .write_en(w_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) w_sh_read0_0 (
        .clk(w_sh_read0_0_clk),
        .done(w_sh_read0_0_done),
        .in(w_sh_read0_0_in),
        .out(w_sh_read0_0_out),
        .write_en(w_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) x0 (
        .addr0(x0_addr0),
        .clk(x0_clk),
        .done(x0_done),
        .read_data(x0_read_data),
        .write_data(x0_write_data),
        .write_en(x0_write_en)
    );
    std_reg # (
        .width(32)
    ) x_int_read0_0 (
        .clk(x_int_read0_0_clk),
        .done(x_int_read0_0_done),
        .in(x_int_read0_0_in),
        .out(x_int_read0_0_out),
        .write_en(x_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) x_read0_0 (
        .clk(x_read0_0_clk),
        .done(x_read0_0_done),
        .in(x_read0_0_in),
        .out(x_read0_0_out),
        .write_en(x_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) x_sh_read0_0 (
        .clk(x_sh_read0_0_clk),
        .done(x_sh_read0_0_done),
        .in(x_sh_read0_0_in),
        .out(x_sh_read0_0_out),
        .write_en(x_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) y0 (
        .addr0(y0_addr0),
        .clk(y0_clk),
        .done(y0_done),
        .read_data(y0_read_data),
        .write_data(y0_write_data),
        .write_en(y0_write_en)
    );
    std_reg # (
        .width(32)
    ) y_int_read0_0 (
        .clk(y_int_read0_0_clk),
        .done(y_int_read0_0_done),
        .in(y_int_read0_0_in),
        .out(y_int_read0_0_out),
        .write_en(y_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) y_read0_0 (
        .clk(y_read0_0_clk),
        .done(y_read0_0_done),
        .in(y_read0_0_in),
        .out(y_read0_0_out),
        .write_en(y_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) y_sh_read0_0 (
        .clk(y_sh_read0_0_clk),
        .done(y_sh_read0_0_done),
        .in(y_sh_read0_0_in),
        .out(y_sh_read0_0_out),
        .write_en(y_sh_read0_0_write_en)
    );
    std_mem_d1 # (
        .idx_size(7),
        .size(64),
        .width(32)
    ) z0 (
        .addr0(z0_addr0),
        .clk(z0_clk),
        .done(z0_done),
        .read_data(z0_read_data),
        .write_data(z0_write_data),
        .write_en(z0_write_en)
    );
    std_reg # (
        .width(32)
    ) z_int_read0_0 (
        .clk(z_int_read0_0_clk),
        .done(z_int_read0_0_done),
        .in(z_int_read0_0_in),
        .out(z_int_read0_0_out),
        .write_en(z_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) z_sh_read0_0 (
        .clk(z_sh_read0_0_clk),
        .done(z_sh_read0_0_done),
        .in(z_sh_read0_0_in),
        .out(z_sh_read0_0_out),
        .write_en(z_sh_read0_0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset (
        .clk(par_reset_clk),
        .done(par_reset_done),
        .in(par_reset_in),
        .out(par_reset_out),
        .write_en(par_reset_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg (
        .clk(par_done_reg_clk),
        .done(par_done_reg_done),
        .in(par_done_reg_in),
        .out(par_done_reg_out),
        .write_en(par_done_reg_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg0 (
        .clk(par_done_reg0_clk),
        .done(par_done_reg0_done),
        .in(par_done_reg0_in),
        .out(par_done_reg0_out),
        .write_en(par_done_reg0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset0 (
        .clk(par_reset0_clk),
        .done(par_reset0_done),
        .in(par_reset0_in),
        .out(par_reset0_out),
        .write_en(par_reset0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg1 (
        .clk(par_done_reg1_clk),
        .done(par_done_reg1_done),
        .in(par_done_reg1_in),
        .out(par_done_reg1_out),
        .write_en(par_done_reg1_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg2 (
        .clk(par_done_reg2_clk),
        .done(par_done_reg2_done),
        .in(par_done_reg2_in),
        .out(par_done_reg2_out),
        .write_en(par_done_reg2_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset1 (
        .clk(par_reset1_clk),
        .done(par_reset1_done),
        .in(par_reset1_in),
        .out(par_reset1_out),
        .write_en(par_reset1_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg3 (
        .clk(par_done_reg3_clk),
        .done(par_done_reg3_done),
        .in(par_done_reg3_in),
        .out(par_done_reg3_out),
        .write_en(par_done_reg3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg4 (
        .clk(par_done_reg4_clk),
        .done(par_done_reg4_done),
        .in(par_done_reg4_in),
        .out(par_done_reg4_out),
        .write_en(par_done_reg4_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset2 (
        .clk(par_reset2_clk),
        .done(par_reset2_done),
        .in(par_reset2_in),
        .out(par_reset2_out),
        .write_en(par_reset2_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg5 (
        .clk(par_done_reg5_clk),
        .done(par_done_reg5_done),
        .in(par_done_reg5_in),
        .out(par_done_reg5_out),
        .write_en(par_done_reg5_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg6 (
        .clk(par_done_reg6_clk),
        .done(par_done_reg6_done),
        .in(par_done_reg6_in),
        .out(par_done_reg6_out),
        .write_en(par_done_reg6_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset3 (
        .clk(par_reset3_clk),
        .done(par_reset3_done),
        .in(par_reset3_in),
        .out(par_reset3_out),
        .write_en(par_reset3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg7 (
        .clk(par_done_reg7_clk),
        .done(par_done_reg7_done),
        .in(par_done_reg7_in),
        .out(par_done_reg7_out),
        .write_en(par_done_reg7_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg8 (
        .clk(par_done_reg8_clk),
        .done(par_done_reg8_done),
        .in(par_done_reg8_in),
        .out(par_done_reg8_out),
        .write_en(par_done_reg8_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset4 (
        .clk(par_reset4_clk),
        .done(par_reset4_done),
        .in(par_reset4_in),
        .out(par_reset4_out),
        .write_en(par_reset4_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg9 (
        .clk(par_done_reg9_clk),
        .done(par_done_reg9_done),
        .in(par_done_reg9_in),
        .out(par_done_reg9_out),
        .write_en(par_done_reg9_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg10 (
        .clk(par_done_reg10_clk),
        .done(par_done_reg10_done),
        .in(par_done_reg10_in),
        .out(par_done_reg10_out),
        .write_en(par_done_reg10_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset5 (
        .clk(par_reset5_clk),
        .done(par_reset5_done),
        .in(par_reset5_in),
        .out(par_reset5_out),
        .write_en(par_reset5_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg11 (
        .clk(par_done_reg11_clk),
        .done(par_done_reg11_done),
        .in(par_done_reg11_in),
        .out(par_done_reg11_out),
        .write_en(par_done_reg11_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg12 (
        .clk(par_done_reg12_clk),
        .done(par_done_reg12_done),
        .in(par_done_reg12_in),
        .out(par_done_reg12_out),
        .write_en(par_done_reg12_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .write_en(fsm_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed (
        .clk(cond_computed_clk),
        .done(cond_computed_done),
        .in(cond_computed_in),
        .out(cond_computed_out),
        .write_en(cond_computed_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored (
        .clk(cond_stored_clk),
        .done(cond_stored_done),
        .in(cond_stored_in),
        .out(cond_stored_out),
        .write_en(cond_stored_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg (
        .clk(done_reg_clk),
        .done(done_reg_done),
        .in(done_reg_in),
        .out(done_reg_out),
        .write_en(done_reg_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm0 (
        .clk(fsm0_clk),
        .done(fsm0_done),
        .in(fsm0_in),
        .out(fsm0_out),
        .write_en(fsm0_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm1 (
        .clk(fsm1_clk),
        .done(fsm1_done),
        .in(fsm1_in),
        .out(fsm1_out),
        .write_en(fsm1_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed0 (
        .clk(cond_computed0_clk),
        .done(cond_computed0_done),
        .in(cond_computed0_in),
        .out(cond_computed0_out),
        .write_en(cond_computed0_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored0 (
        .clk(cond_stored0_clk),
        .done(cond_stored0_done),
        .in(cond_stored0_in),
        .out(cond_stored0_out),
        .write_en(cond_stored0_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg0 (
        .clk(done_reg0_clk),
        .done(done_reg0_done),
        .in(done_reg0_in),
        .out(done_reg0_out),
        .write_en(done_reg0_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm2 (
        .clk(fsm2_clk),
        .done(fsm2_done),
        .in(fsm2_in),
        .out(fsm2_out),
        .write_en(fsm2_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed1 (
        .clk(cond_computed1_clk),
        .done(cond_computed1_done),
        .in(cond_computed1_in),
        .out(cond_computed1_out),
        .write_en(cond_computed1_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored1 (
        .clk(cond_stored1_clk),
        .done(cond_stored1_done),
        .in(cond_stored1_in),
        .out(cond_stored1_out),
        .write_en(cond_stored1_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg1 (
        .clk(done_reg1_clk),
        .done(done_reg1_done),
        .in(done_reg1_in),
        .out(done_reg1_out),
        .write_en(done_reg1_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm3 (
        .clk(fsm3_clk),
        .done(fsm3_done),
        .in(fsm3_in),
        .out(fsm3_out),
        .write_en(fsm3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset6 (
        .clk(par_reset6_clk),
        .done(par_reset6_done),
        .in(par_reset6_in),
        .out(par_reset6_out),
        .write_en(par_reset6_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg13 (
        .clk(par_done_reg13_clk),
        .done(par_done_reg13_done),
        .in(par_done_reg13_in),
        .out(par_done_reg13_out),
        .write_en(par_done_reg13_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg14 (
        .clk(par_done_reg14_clk),
        .done(par_done_reg14_done),
        .in(par_done_reg14_in),
        .out(par_done_reg14_out),
        .write_en(par_done_reg14_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg15 (
        .clk(par_done_reg15_clk),
        .done(par_done_reg15_done),
        .in(par_done_reg15_in),
        .out(par_done_reg15_out),
        .write_en(par_done_reg15_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg16 (
        .clk(par_done_reg16_clk),
        .done(par_done_reg16_done),
        .in(par_done_reg16_in),
        .out(par_done_reg16_out),
        .write_en(par_done_reg16_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset7 (
        .clk(par_reset7_clk),
        .done(par_reset7_done),
        .in(par_reset7_in),
        .out(par_reset7_out),
        .write_en(par_reset7_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg17 (
        .clk(par_done_reg17_clk),
        .done(par_done_reg17_done),
        .in(par_done_reg17_in),
        .out(par_done_reg17_out),
        .write_en(par_done_reg17_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg18 (
        .clk(par_done_reg18_clk),
        .done(par_done_reg18_done),
        .in(par_done_reg18_in),
        .out(par_done_reg18_out),
        .write_en(par_done_reg18_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg19 (
        .clk(par_done_reg19_clk),
        .done(par_done_reg19_done),
        .in(par_done_reg19_in),
        .out(par_done_reg19_out),
        .write_en(par_done_reg19_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg20 (
        .clk(par_done_reg20_clk),
        .done(par_done_reg20_done),
        .in(par_done_reg20_in),
        .out(par_done_reg20_out),
        .write_en(par_done_reg20_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm4 (
        .clk(fsm4_clk),
        .done(fsm4_done),
        .in(fsm4_in),
        .out(fsm4_out),
        .write_en(fsm4_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset8 (
        .clk(par_reset8_clk),
        .done(par_reset8_done),
        .in(par_reset8_in),
        .out(par_reset8_out),
        .write_en(par_reset8_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg21 (
        .clk(par_done_reg21_clk),
        .done(par_done_reg21_done),
        .in(par_done_reg21_in),
        .out(par_done_reg21_out),
        .write_en(par_done_reg21_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg22 (
        .clk(par_done_reg22_clk),
        .done(par_done_reg22_done),
        .in(par_done_reg22_in),
        .out(par_done_reg22_out),
        .write_en(par_done_reg22_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm5 (
        .clk(fsm5_clk),
        .done(fsm5_done),
        .in(fsm5_in),
        .out(fsm5_out),
        .write_en(fsm5_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed2 (
        .clk(cond_computed2_clk),
        .done(cond_computed2_done),
        .in(cond_computed2_in),
        .out(cond_computed2_out),
        .write_en(cond_computed2_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored2 (
        .clk(cond_stored2_clk),
        .done(cond_stored2_done),
        .in(cond_stored2_in),
        .out(cond_stored2_out),
        .write_en(cond_stored2_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg2 (
        .clk(done_reg2_clk),
        .done(done_reg2_done),
        .in(done_reg2_in),
        .out(done_reg2_out),
        .write_en(done_reg2_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm6 (
        .clk(fsm6_clk),
        .done(fsm6_done),
        .in(fsm6_in),
        .out(fsm6_out),
        .write_en(fsm6_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed3 (
        .clk(cond_computed3_clk),
        .done(cond_computed3_done),
        .in(cond_computed3_in),
        .out(cond_computed3_out),
        .write_en(cond_computed3_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored3 (
        .clk(cond_stored3_clk),
        .done(cond_stored3_done),
        .in(cond_stored3_in),
        .out(cond_stored3_out),
        .write_en(cond_stored3_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg3 (
        .clk(done_reg3_clk),
        .done(done_reg3_done),
        .in(done_reg3_in),
        .out(done_reg3_out),
        .write_en(done_reg3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset9 (
        .clk(par_reset9_clk),
        .done(par_reset9_done),
        .in(par_reset9_in),
        .out(par_reset9_out),
        .write_en(par_reset9_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg23 (
        .clk(par_done_reg23_clk),
        .done(par_done_reg23_done),
        .in(par_done_reg23_in),
        .out(par_done_reg23_out),
        .write_en(par_done_reg23_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg24 (
        .clk(par_done_reg24_clk),
        .done(par_done_reg24_done),
        .in(par_done_reg24_in),
        .out(par_done_reg24_out),
        .write_en(par_done_reg24_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm7 (
        .clk(fsm7_clk),
        .done(fsm7_done),
        .in(fsm7_in),
        .out(fsm7_out),
        .write_en(fsm7_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed4 (
        .clk(cond_computed4_clk),
        .done(cond_computed4_done),
        .in(cond_computed4_in),
        .out(cond_computed4_out),
        .write_en(cond_computed4_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored4 (
        .clk(cond_stored4_clk),
        .done(cond_stored4_done),
        .in(cond_stored4_in),
        .out(cond_stored4_out),
        .write_en(cond_stored4_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg4 (
        .clk(done_reg4_clk),
        .done(done_reg4_done),
        .in(done_reg4_in),
        .out(done_reg4_out),
        .write_en(done_reg4_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm8 (
        .clk(fsm8_clk),
        .done(fsm8_done),
        .in(fsm8_in),
        .out(fsm8_out),
        .write_en(fsm8_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed5 (
        .clk(cond_computed5_clk),
        .done(cond_computed5_done),
        .in(cond_computed5_in),
        .out(cond_computed5_out),
        .write_en(cond_computed5_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored5 (
        .clk(cond_stored5_clk),
        .done(cond_stored5_done),
        .in(cond_stored5_in),
        .out(cond_stored5_out),
        .write_en(cond_stored5_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg5 (
        .clk(done_reg5_clk),
        .done(done_reg5_done),
        .in(done_reg5_in),
        .out(done_reg5_out),
        .write_en(done_reg5_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset10 (
        .clk(par_reset10_clk),
        .done(par_reset10_done),
        .in(par_reset10_in),
        .out(par_reset10_out),
        .write_en(par_reset10_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg25 (
        .clk(par_done_reg25_clk),
        .done(par_done_reg25_done),
        .in(par_done_reg25_in),
        .out(par_done_reg25_out),
        .write_en(par_done_reg25_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg26 (
        .clk(par_done_reg26_clk),
        .done(par_done_reg26_done),
        .in(par_done_reg26_in),
        .out(par_done_reg26_out),
        .write_en(par_done_reg26_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm9 (
        .clk(fsm9_clk),
        .done(fsm9_done),
        .in(fsm9_in),
        .out(fsm9_out),
        .write_en(fsm9_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed6 (
        .clk(cond_computed6_clk),
        .done(cond_computed6_done),
        .in(cond_computed6_in),
        .out(cond_computed6_out),
        .write_en(cond_computed6_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored6 (
        .clk(cond_stored6_clk),
        .done(cond_stored6_done),
        .in(cond_stored6_in),
        .out(cond_stored6_out),
        .write_en(cond_stored6_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg6 (
        .clk(done_reg6_clk),
        .done(done_reg6_done),
        .in(done_reg6_in),
        .out(done_reg6_out),
        .write_en(done_reg6_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset11 (
        .clk(par_reset11_clk),
        .done(par_reset11_done),
        .in(par_reset11_in),
        .out(par_reset11_out),
        .write_en(par_reset11_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg27 (
        .clk(par_done_reg27_clk),
        .done(par_done_reg27_done),
        .in(par_done_reg27_in),
        .out(par_done_reg27_out),
        .write_en(par_done_reg27_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg28 (
        .clk(par_done_reg28_clk),
        .done(par_done_reg28_done),
        .in(par_done_reg28_in),
        .out(par_done_reg28_out),
        .write_en(par_done_reg28_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm10 (
        .clk(fsm10_clk),
        .done(fsm10_done),
        .in(fsm10_in),
        .out(fsm10_out),
        .write_en(fsm10_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed7 (
        .clk(cond_computed7_clk),
        .done(cond_computed7_done),
        .in(cond_computed7_in),
        .out(cond_computed7_out),
        .write_en(cond_computed7_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored7 (
        .clk(cond_stored7_clk),
        .done(cond_stored7_done),
        .in(cond_stored7_in),
        .out(cond_stored7_out),
        .write_en(cond_stored7_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg7 (
        .clk(done_reg7_clk),
        .done(done_reg7_done),
        .in(done_reg7_in),
        .out(done_reg7_out),
        .write_en(done_reg7_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm11 (
        .clk(fsm11_clk),
        .done(fsm11_done),
        .in(fsm11_in),
        .out(fsm11_out),
        .write_en(fsm11_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed8 (
        .clk(cond_computed8_clk),
        .done(cond_computed8_done),
        .in(cond_computed8_in),
        .out(cond_computed8_out),
        .write_en(cond_computed8_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored8 (
        .clk(cond_stored8_clk),
        .done(cond_stored8_done),
        .in(cond_stored8_in),
        .out(cond_stored8_out),
        .write_en(cond_stored8_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg8 (
        .clk(done_reg8_clk),
        .done(done_reg8_done),
        .in(done_reg8_in),
        .out(done_reg8_out),
        .write_en(done_reg8_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset12 (
        .clk(par_reset12_clk),
        .done(par_reset12_done),
        .in(par_reset12_in),
        .out(par_reset12_out),
        .write_en(par_reset12_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg29 (
        .clk(par_done_reg29_clk),
        .done(par_done_reg29_done),
        .in(par_done_reg29_in),
        .out(par_done_reg29_out),
        .write_en(par_done_reg29_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg30 (
        .clk(par_done_reg30_clk),
        .done(par_done_reg30_done),
        .in(par_done_reg30_in),
        .out(par_done_reg30_out),
        .write_en(par_done_reg30_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset13 (
        .clk(par_reset13_clk),
        .done(par_reset13_done),
        .in(par_reset13_in),
        .out(par_reset13_out),
        .write_en(par_reset13_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg31 (
        .clk(par_done_reg31_clk),
        .done(par_done_reg31_done),
        .in(par_done_reg31_in),
        .out(par_done_reg31_out),
        .write_en(par_done_reg31_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg32 (
        .clk(par_done_reg32_clk),
        .done(par_done_reg32_done),
        .in(par_done_reg32_in),
        .out(par_done_reg32_out),
        .write_en(par_done_reg32_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset14 (
        .clk(par_reset14_clk),
        .done(par_reset14_done),
        .in(par_reset14_in),
        .out(par_reset14_out),
        .write_en(par_reset14_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg33 (
        .clk(par_done_reg33_clk),
        .done(par_done_reg33_done),
        .in(par_done_reg33_in),
        .out(par_done_reg33_out),
        .write_en(par_done_reg33_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg34 (
        .clk(par_done_reg34_clk),
        .done(par_done_reg34_done),
        .in(par_done_reg34_in),
        .out(par_done_reg34_out),
        .write_en(par_done_reg34_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset15 (
        .clk(par_reset15_clk),
        .done(par_reset15_done),
        .in(par_reset15_in),
        .out(par_reset15_out),
        .write_en(par_reset15_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg35 (
        .clk(par_done_reg35_clk),
        .done(par_done_reg35_done),
        .in(par_done_reg35_in),
        .out(par_done_reg35_out),
        .write_en(par_done_reg35_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg36 (
        .clk(par_done_reg36_clk),
        .done(par_done_reg36_done),
        .in(par_done_reg36_in),
        .out(par_done_reg36_out),
        .write_en(par_done_reg36_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset16 (
        .clk(par_reset16_clk),
        .done(par_reset16_done),
        .in(par_reset16_in),
        .out(par_reset16_out),
        .write_en(par_reset16_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg37 (
        .clk(par_done_reg37_clk),
        .done(par_done_reg37_done),
        .in(par_done_reg37_in),
        .out(par_done_reg37_out),
        .write_en(par_done_reg37_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg38 (
        .clk(par_done_reg38_clk),
        .done(par_done_reg38_done),
        .in(par_done_reg38_in),
        .out(par_done_reg38_out),
        .write_en(par_done_reg38_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset17 (
        .clk(par_reset17_clk),
        .done(par_reset17_done),
        .in(par_reset17_in),
        .out(par_reset17_out),
        .write_en(par_reset17_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg39 (
        .clk(par_done_reg39_clk),
        .done(par_done_reg39_done),
        .in(par_done_reg39_in),
        .out(par_done_reg39_out),
        .write_en(par_done_reg39_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg40 (
        .clk(par_done_reg40_clk),
        .done(par_done_reg40_done),
        .in(par_done_reg40_in),
        .out(par_done_reg40_out),
        .write_en(par_done_reg40_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset18 (
        .clk(par_reset18_clk),
        .done(par_reset18_done),
        .in(par_reset18_in),
        .out(par_reset18_out),
        .write_en(par_reset18_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg41 (
        .clk(par_done_reg41_clk),
        .done(par_done_reg41_done),
        .in(par_done_reg41_in),
        .out(par_done_reg41_out),
        .write_en(par_done_reg41_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg42 (
        .clk(par_done_reg42_clk),
        .done(par_done_reg42_done),
        .in(par_done_reg42_in),
        .out(par_done_reg42_out),
        .write_en(par_done_reg42_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm12 (
        .clk(fsm12_clk),
        .done(fsm12_done),
        .in(fsm12_in),
        .out(fsm12_out),
        .write_en(fsm12_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed9 (
        .clk(cond_computed9_clk),
        .done(cond_computed9_done),
        .in(cond_computed9_in),
        .out(cond_computed9_out),
        .write_en(cond_computed9_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored9 (
        .clk(cond_stored9_clk),
        .done(cond_stored9_done),
        .in(cond_stored9_in),
        .out(cond_stored9_out),
        .write_en(cond_stored9_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg9 (
        .clk(done_reg9_clk),
        .done(done_reg9_done),
        .in(done_reg9_in),
        .out(done_reg9_out),
        .write_en(done_reg9_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm13 (
        .clk(fsm13_clk),
        .done(fsm13_done),
        .in(fsm13_in),
        .out(fsm13_out),
        .write_en(fsm13_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm14 (
        .clk(fsm14_clk),
        .done(fsm14_done),
        .in(fsm14_in),
        .out(fsm14_out),
        .write_en(fsm14_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed10 (
        .clk(cond_computed10_clk),
        .done(cond_computed10_done),
        .in(cond_computed10_in),
        .out(cond_computed10_out),
        .write_en(cond_computed10_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored10 (
        .clk(cond_stored10_clk),
        .done(cond_stored10_done),
        .in(cond_stored10_in),
        .out(cond_stored10_out),
        .write_en(cond_stored10_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg10 (
        .clk(done_reg10_clk),
        .done(done_reg10_done),
        .in(done_reg10_in),
        .out(done_reg10_out),
        .write_en(done_reg10_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm15 (
        .clk(fsm15_clk),
        .done(fsm15_done),
        .in(fsm15_in),
        .out(fsm15_out),
        .write_en(fsm15_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed11 (
        .clk(cond_computed11_clk),
        .done(cond_computed11_done),
        .in(cond_computed11_in),
        .out(cond_computed11_out),
        .write_en(cond_computed11_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored11 (
        .clk(cond_stored11_clk),
        .done(cond_stored11_done),
        .in(cond_stored11_in),
        .out(cond_stored11_out),
        .write_en(cond_stored11_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg11 (
        .clk(done_reg11_clk),
        .done(done_reg11_done),
        .in(done_reg11_in),
        .out(done_reg11_out),
        .write_en(done_reg11_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm16 (
        .clk(fsm16_clk),
        .done(fsm16_done),
        .in(fsm16_in),
        .out(fsm16_out),
        .write_en(fsm16_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset19 (
        .clk(par_reset19_clk),
        .done(par_reset19_done),
        .in(par_reset19_in),
        .out(par_reset19_out),
        .write_en(par_reset19_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg43 (
        .clk(par_done_reg43_clk),
        .done(par_done_reg43_done),
        .in(par_done_reg43_in),
        .out(par_done_reg43_out),
        .write_en(par_done_reg43_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg44 (
        .clk(par_done_reg44_clk),
        .done(par_done_reg44_done),
        .in(par_done_reg44_in),
        .out(par_done_reg44_out),
        .write_en(par_done_reg44_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm17 (
        .clk(fsm17_clk),
        .done(fsm17_done),
        .in(fsm17_in),
        .out(fsm17_out),
        .write_en(fsm17_write_en)
    );
    always_comb begin
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A0_0_addr0 = rsh1_out;
        end else if((~(par_done_reg22_out | old_0_done) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            A0_0_addr0 = i2_out;
        end else if((((fsm5_out == 32'd2) & ~A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            A0_0_addr0 = i2_out;
        end else if((~(par_done_reg23_out | A_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            A0_0_addr0 = j2_out;
        end else if((~(par_done_reg27_out | A_read1_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            A0_0_addr0 = i5_out;
        end else if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A0_0_addr0 = rsh1_out;
        end else A0_0_addr0 = 7'd0;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A0_0_addr1 = rsh0_out;
        end else if((~(par_done_reg22_out | old_0_done) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            A0_0_addr1 = j1_out;
        end else if((((fsm5_out == 32'd2) & ~A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            A0_0_addr1 = j1_out;
        end else if((~(par_done_reg23_out | A_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            A0_0_addr1 = i3_out;
        end else if((~(par_done_reg27_out | A_read1_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            A0_0_addr1 = j3_out;
        end else if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A0_0_addr1 = rsh0_out;
        end else A0_0_addr1 = 7'd0;
        A0_0_clk = clk;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A0_0_write_data = A_int_read0_0_out;
        end else if((((fsm5_out == 32'd2) & ~A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            A0_0_write_data = add10_out;
        end else A0_0_write_data = 32'd0;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A0_0_write_en = 1'd1;
        end else if((((fsm5_out == 32'd2) & ~A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            A0_0_write_en = 1'd1;
        end else A0_0_write_en = 1'd0;
        A_int_read0_0_clk = clk;
        if((((fsm1_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A_int_read0_0_in = A_int0_0_read_data;
        end else A_int_read0_0_in = 32'd0;
        if((((fsm1_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A_int_read0_0_write_en = 1'd1;
        end else A_int_read0_0_write_en = 1'd0;
        A_read0_0_clk = clk;
        if((~(par_done_reg23_out | A_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            A_read0_0_in = A0_0_read_data;
        end else A_read0_0_in = 32'd0;
        if((~(par_done_reg23_out | A_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            A_read0_0_write_en = 1'd1;
        end else A_read0_0_write_en = 1'd0;
        A_read1_0_clk = clk;
        if((~(par_done_reg27_out | A_read1_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            A_read1_0_in = A0_0_read_data;
        end else A_read1_0_in = 32'd0;
        if((~(par_done_reg27_out | A_read1_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            A_read1_0_write_en = 1'd1;
        end else A_read1_0_write_en = 1'd0;
        A_sh_read0_0_clk = clk;
        if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A_sh_read0_0_in = A0_0_read_data;
        end else A_sh_read0_0_in = 32'd0;
        if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A_sh_read0_0_write_en = 1'd1;
        end else A_sh_read0_0_write_en = 1'd0;
        if((((fsm1_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A_int0_0_addr0 = i1_out;
        end else if((((fsm14_out == 32'd1) & ~A_int0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A_int0_0_addr0 = i7_out;
        end else A_int0_0_addr0 = 7'd0;
        if((((fsm1_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            A_int0_0_addr1 = j0_out;
        end else if((((fsm14_out == 32'd1) & ~A_int0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A_int0_0_addr1 = j4_out;
        end else A_int0_0_addr1 = 7'd0;
        A_int0_0_clk = clk;
        if((((fsm14_out == 32'd1) & ~A_int0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A_int0_0_write_data = A_sh_read0_0_out;
        end else A_int0_0_write_data = 32'd0;
        if((((fsm14_out == 32'd1) & ~A_int0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            A_int0_0_write_en = 1'd1;
        end else A_int0_0_write_en = 1'd0;
        if((~(par_done_reg13_out | alpha__0_done) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            alpha_int0_addr0 = const0_out;
        end else alpha_int0_addr0 = 1'd0;
        alpha_int0_clk = clk;
        if((~(par_done_reg14_out | beta__0_done) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            beta_int0_addr0 = const1_out;
        end else beta_int0_addr0 = 1'd0;
        beta_int0_clk = clk;
        if((fsm17_out == 32'd10)) begin
            done = 1'd1;
        end else if((fsm17_out == 32'd10)) begin
            done = 1'd1;
        end else done = 1'd0;
        if((((fsm_out == 32'd0) & ~u1_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            u1_int0_addr0 = i0_out;
        end else if((~(par_done_reg29_out | u1_int0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u1_int0_addr0 = i6_out;
        end else u1_int0_addr0 = 7'd0;
        u1_int0_clk = clk;
        if((~(par_done_reg29_out | u1_int0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u1_int0_write_data = u1_sh_read0_0_out;
        end else u1_int0_write_data = 32'd0;
        if((~(par_done_reg29_out | u1_int0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u1_int0_write_en = 1'd1;
        end else u1_int0_write_en = 1'd0;
        if((~(par_done_reg33_out | u2_int0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u2_int0_addr0 = i6_out;
        end else if((~(par_done_reg2_out | u2_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u2_int0_addr0 = i0_out;
        end else u2_int0_addr0 = 7'd0;
        u2_int0_clk = clk;
        if((~(par_done_reg33_out | u2_int0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u2_int0_write_data = u2_sh_read0_0_out;
        end else u2_int0_write_data = 32'd0;
        if((~(par_done_reg33_out | u2_int0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u2_int0_write_en = 1'd1;
        end else u2_int0_write_en = 1'd0;
        if((~(par_done_reg0_out | v1_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v1_int0_addr0 = i0_out;
        end else if((~(par_done_reg31_out | v1_int0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v1_int0_addr0 = i6_out;
        end else v1_int0_addr0 = 7'd0;
        v1_int0_clk = clk;
        if((~(par_done_reg31_out | v1_int0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v1_int0_write_data = v1_sh_read0_0_out;
        end else v1_int0_write_data = 32'd0;
        if((~(par_done_reg31_out | v1_int0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v1_int0_write_en = 1'd1;
        end else v1_int0_write_en = 1'd0;
        if((~(par_done_reg35_out | v2_int0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v2_int0_addr0 = i6_out;
        end else if((~(par_done_reg4_out | v2_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v2_int0_addr0 = i0_out;
        end else v2_int0_addr0 = 7'd0;
        v2_int0_clk = clk;
        if((~(par_done_reg35_out | v2_int0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v2_int0_write_data = v2_sh_read0_0_out;
        end else v2_int0_write_data = 32'd0;
        if((~(par_done_reg35_out | v2_int0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v2_int0_write_en = 1'd1;
        end else v2_int0_write_en = 1'd0;
        if((~(par_done_reg6_out | w_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            w_int0_addr0 = i0_out;
        end else if((~(par_done_reg37_out | w_int0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            w_int0_addr0 = i6_out;
        end else w_int0_addr0 = 7'd0;
        w_int0_clk = clk;
        if((~(par_done_reg37_out | w_int0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            w_int0_write_data = w_sh_read0_0_out;
        end else w_int0_write_data = 32'd0;
        if((~(par_done_reg37_out | w_int0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            w_int0_write_en = 1'd1;
        end else w_int0_write_en = 1'd0;
        if((~(par_done_reg8_out | x_int_read0_0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            x_int0_addr0 = i0_out;
        end else if((~(par_done_reg39_out | x_int0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            x_int0_addr0 = i6_out;
        end else x_int0_addr0 = 7'd0;
        x_int0_clk = clk;
        if((~(par_done_reg39_out | x_int0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            x_int0_write_data = x_sh_read0_0_out;
        end else x_int0_write_data = 32'd0;
        if((~(par_done_reg39_out | x_int0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            x_int0_write_en = 1'd1;
        end else x_int0_write_en = 1'd0;
        if((~(par_done_reg10_out | y_int_read0_0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            y_int0_addr0 = i0_out;
        end else if((~(par_done_reg41_out | y_int0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            y_int0_addr0 = i6_out;
        end else y_int0_addr0 = 7'd0;
        y_int0_clk = clk;
        if((~(par_done_reg41_out | y_int0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            y_int0_write_data = y_sh_read0_0_out;
        end else y_int0_write_data = 32'd0;
        if((~(par_done_reg41_out | y_int0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            y_int0_write_en = 1'd1;
        end else y_int0_write_en = 1'd0;
        if((~(par_done_reg12_out | z_int_read0_0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            z_int0_addr0 = i0_out;
        end else if((((fsm12_out == 32'd8) & ~z_int0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            z_int0_addr0 = i6_out;
        end else z_int0_addr0 = 7'd0;
        z_int0_clk = clk;
        if((((fsm12_out == 32'd8) & ~z_int0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            z_int0_write_data = z_sh_read0_0_out;
        end else z_int0_write_data = 32'd0;
        if((((fsm12_out == 32'd8) & ~z_int0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            z_int0_write_en = 1'd1;
        end else z_int0_write_en = 1'd0;
        if((((fsm1_out == 32'd2) & ~j0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            add0_left = j0_out;
        end else if((((fsm2_out == 32'd2) & ~i1_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            add0_left = i1_out;
        end else if((((fsm5_out == 32'd3) & ~j1_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            add0_left = j1_out;
        end else if((((fsm6_out == 32'd2) & ~i2_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            add0_left = i2_out;
        end else if((((fsm7_out == 32'd5) & ~j2_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            add0_left = j2_out;
        end else if((((fsm8_out == 32'd2) & ~i3_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            add0_left = i3_out;
        end else if((((fsm9_out == 32'd2) & ~i4_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            add0_left = i4_out;
        end else if((((fsm10_out == 32'd5) & ~j3_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            add0_left = j3_out;
        end else if((((fsm11_out == 32'd2) & ~i5_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            add0_left = i5_out;
        end else if((((fsm14_out == 32'd2) & ~j4_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            add0_left = j4_out;
        end else if((((fsm15_out == 32'd2) & ~i7_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            add0_left = i7_out;
        end else add0_left = 7'd0;
        if((((fsm1_out == 32'd2) & ~j0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            add0_right = const12_out;
        end else if((((fsm2_out == 32'd2) & ~i1_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            add0_right = const12_out;
        end else if((((fsm5_out == 32'd3) & ~j1_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            add0_right = const12_out;
        end else if((((fsm6_out == 32'd2) & ~i2_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            add0_right = const12_out;
        end else if((((fsm7_out == 32'd5) & ~j2_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            add0_right = const12_out;
        end else if((((fsm8_out == 32'd2) & ~i3_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            add0_right = const12_out;
        end else if((((fsm9_out == 32'd2) & ~i4_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            add0_right = const12_out;
        end else if((((fsm10_out == 32'd5) & ~j3_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            add0_right = const12_out;
        end else if((((fsm11_out == 32'd2) & ~i5_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            add0_right = const12_out;
        end else if((((fsm14_out == 32'd2) & ~j4_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            add0_right = const12_out;
        end else if((((fsm15_out == 32'd2) & ~i7_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            add0_right = const12_out;
        end else add0_right = 7'd0;
        if((((fsm_out == 32'd9) & ~i0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            add1_left = i0_out;
        end else if((((fsm12_out == 32'd9) & ~i6_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            add1_left = i6_out;
        end else add1_left = 7'd0;
        if((((fsm_out == 32'd9) & ~i0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            add1_right = const19_out;
        end else if((((fsm12_out == 32'd9) & ~i6_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            add1_right = const19_out;
        end else add1_right = 7'd0;
        if((((fsm4_out == 32'd2) & ~tmp1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            add10_left = bin_read0_0_out;
        end else if((((fsm5_out == 32'd2) & ~A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            add10_left = old_0_out;
        end else if((((fsm7_out == 32'd4) & ~x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            add10_left = x0_read_data;
        end else if((((fsm9_out == 32'd1) & ~x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            add10_left = old_1_out;
        end else if((((fsm10_out == 32'd4) & ~w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            add10_left = w0_read_data;
        end else add10_left = 32'd0;
        if((((fsm4_out == 32'd2) & ~tmp1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            add10_right = bin_read1_0_out;
        end else if((((fsm5_out == 32'd2) & ~A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            add10_right = tmp1_0_out;
        end else if((((fsm7_out == 32'd4) & ~x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            add10_right = tmp2_0_out;
        end else if((((fsm9_out == 32'd1) & ~x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            add10_right = tmp3_0_out;
        end else if((((fsm10_out == 32'd4) & ~w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            add10_right = tmp4_0_out;
        end else add10_right = 32'd0;
        alpha__0_clk = clk;
        if((~(par_done_reg13_out | alpha__0_done) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            alpha__0_in = alpha_int0_read_data;
        end else alpha__0_in = 32'd0;
        if((~(par_done_reg13_out | alpha__0_done) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            alpha__0_write_en = 1'd1;
        end else alpha__0_write_en = 1'd0;
        beta__0_clk = clk;
        if((~(par_done_reg14_out | beta__0_done) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            beta__0_in = beta_int0_read_data;
        end else beta__0_in = 32'd0;
        if((~(par_done_reg14_out | beta__0_done) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            beta__0_write_en = 1'd1;
        end else beta__0_write_en = 1'd0;
        bin_read0_0_clk = clk;
        if((((fsm4_out == 32'd0) & ~bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read0_0_in = mult_pipe0_out;
        end else bin_read0_0_in = 32'd0;
        if((((fsm4_out == 32'd0) & ~bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read0_0_write_en = mult_pipe0_done;
        end else bin_read0_0_write_en = 1'd0;
        bin_read1_0_clk = clk;
        if((((fsm4_out == 32'd1) & ~bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read1_0_in = mult_pipe1_out;
        end else bin_read1_0_in = 32'd0;
        if((((fsm4_out == 32'd1) & ~bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read1_0_write_en = mult_pipe1_done;
        end else bin_read1_0_write_en = 1'd0;
        bin_read2_0_clk = clk;
        if((((fsm7_out == 32'd1) & ~bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            bin_read2_0_in = mult_pipe2_out;
        end else bin_read2_0_in = 32'd0;
        if((((fsm7_out == 32'd1) & ~bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            bin_read2_0_write_en = mult_pipe2_done;
        end else bin_read2_0_write_en = 1'd0;
        bin_read3_0_clk = clk;
        if((((fsm7_out == 32'd2) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            bin_read3_0_in = mult_pipe3_out;
        end else bin_read3_0_in = 32'd0;
        if((((fsm7_out == 32'd2) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            bin_read3_0_write_en = mult_pipe3_done;
        end else bin_read3_0_write_en = 1'd0;
        bin_read4_0_clk = clk;
        if((((fsm10_out == 32'd1) & ~bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            bin_read4_0_in = mult_pipe4_out;
        end else bin_read4_0_in = 32'd0;
        if((((fsm10_out == 32'd1) & ~bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            bin_read4_0_write_en = mult_pipe4_done;
        end else bin_read4_0_write_en = 1'd0;
        bin_read5_0_clk = clk;
        if((((fsm10_out == 32'd2) & ~bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            bin_read5_0_in = mult_pipe5_out;
        end else bin_read5_0_in = 32'd0;
        if((((fsm10_out == 32'd2) & ~bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            bin_read5_0_write_en = mult_pipe5_done;
        end else bin_read5_0_write_en = 1'd0;
        cond_computed_clk = clk;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed_in = 1'd1;
        end else if((((cond_stored_out & cond_computed_out) & (fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed_in = 1'd0;
        end else if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed_in = 1'd0;
        end else cond_computed_in = 1'd0;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed_write_en = 1'd1;
        end else if((((cond_stored_out & cond_computed_out) & (fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed_write_en = 1'd1;
        end else if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed_write_en = 1'd1;
        end else cond_computed_write_en = 1'd0;
        cond_computed0_clk = clk;
        if((((~cond_computed0_out & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_computed0_in = 1'd1;
        end else if((((cond_stored0_out & cond_computed0_out) & (fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_computed0_in = 1'd0;
        end else if(((cond_computed0_out & ~cond_stored0_out) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_computed0_in = 1'd0;
        end else cond_computed0_in = 1'd0;
        if((((~cond_computed0_out & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_computed0_write_en = 1'd1;
        end else if((((cond_stored0_out & cond_computed0_out) & (fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_computed0_write_en = 1'd1;
        end else if(((cond_computed0_out & ~cond_stored0_out) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_computed0_write_en = 1'd1;
        end else cond_computed0_write_en = 1'd0;
        cond_computed1_clk = clk;
        if((((~cond_computed1_out & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed1_in = 1'd1;
        end else if((((cond_stored1_out & cond_computed1_out) & (fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed1_in = 1'd0;
        end else if(((cond_computed1_out & ~cond_stored1_out) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed1_in = 1'd0;
        end else cond_computed1_in = 1'd0;
        if((((~cond_computed1_out & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed1_write_en = 1'd1;
        end else if((((cond_stored1_out & cond_computed1_out) & (fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed1_write_en = 1'd1;
        end else if(((cond_computed1_out & ~cond_stored1_out) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_computed1_write_en = 1'd1;
        end else cond_computed1_write_en = 1'd0;
        cond_computed10_clk = clk;
        if((((~cond_computed10_out & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) & 1'b1) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_computed10_in = 1'd1;
        end else if((((cond_stored10_out & cond_computed10_out) & (fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_computed10_in = 1'd0;
        end else if(((cond_computed10_out & ~cond_stored10_out) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_computed10_in = 1'd0;
        end else cond_computed10_in = 1'd0;
        if((((~cond_computed10_out & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) & 1'b1) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_computed10_write_en = 1'd1;
        end else if((((cond_stored10_out & cond_computed10_out) & (fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_computed10_write_en = 1'd1;
        end else if(((cond_computed10_out & ~cond_stored10_out) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_computed10_write_en = 1'd1;
        end else cond_computed10_write_en = 1'd0;
        cond_computed11_clk = clk;
        if((((~cond_computed11_out & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed11_in = 1'd1;
        end else if((((cond_stored11_out & cond_computed11_out) & (fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed11_in = 1'd0;
        end else if(((cond_computed11_out & ~cond_stored11_out) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed11_in = 1'd0;
        end else cond_computed11_in = 1'd0;
        if((((~cond_computed11_out & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed11_write_en = 1'd1;
        end else if((((cond_stored11_out & cond_computed11_out) & (fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed11_write_en = 1'd1;
        end else if(((cond_computed11_out & ~cond_stored11_out) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed11_write_en = 1'd1;
        end else cond_computed11_write_en = 1'd0;
        cond_computed2_clk = clk;
        if((((~cond_computed2_out & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_in = 1'd1;
        end else if((((cond_stored2_out & cond_computed2_out) & (fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_in = 1'd0;
        end else if(((cond_computed2_out & ~cond_stored2_out) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_in = 1'd0;
        end else cond_computed2_in = 1'd0;
        if((((~cond_computed2_out & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_write_en = 1'd1;
        end else if((((cond_stored2_out & cond_computed2_out) & (fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_write_en = 1'd1;
        end else if(((cond_computed2_out & ~cond_stored2_out) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_write_en = 1'd1;
        end else cond_computed2_write_en = 1'd0;
        cond_computed3_clk = clk;
        if((((~cond_computed3_out & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_in = 1'd1;
        end else if((((cond_stored3_out & cond_computed3_out) & (fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_in = 1'd0;
        end else if(((cond_computed3_out & ~cond_stored3_out) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_in = 1'd0;
        end else cond_computed3_in = 1'd0;
        if((((~cond_computed3_out & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_write_en = 1'd1;
        end else if((((cond_stored3_out & cond_computed3_out) & (fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_write_en = 1'd1;
        end else if(((cond_computed3_out & ~cond_stored3_out) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_write_en = 1'd1;
        end else cond_computed3_write_en = 1'd0;
        cond_computed4_clk = clk;
        if((((~cond_computed4_out & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_computed4_in = 1'd1;
        end else if((((cond_stored4_out & cond_computed4_out) & (fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_computed4_in = 1'd0;
        end else if(((cond_computed4_out & ~cond_stored4_out) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_computed4_in = 1'd0;
        end else cond_computed4_in = 1'd0;
        if((((~cond_computed4_out & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_computed4_write_en = 1'd1;
        end else if((((cond_stored4_out & cond_computed4_out) & (fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_computed4_write_en = 1'd1;
        end else if(((cond_computed4_out & ~cond_stored4_out) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_computed4_write_en = 1'd1;
        end else cond_computed4_write_en = 1'd0;
        cond_computed5_clk = clk;
        if((((~cond_computed5_out & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_computed5_in = 1'd1;
        end else if((((cond_stored5_out & cond_computed5_out) & (fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_computed5_in = 1'd0;
        end else if(((cond_computed5_out & ~cond_stored5_out) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_computed5_in = 1'd0;
        end else cond_computed5_in = 1'd0;
        if((((~cond_computed5_out & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_computed5_write_en = 1'd1;
        end else if((((cond_stored5_out & cond_computed5_out) & (fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_computed5_write_en = 1'd1;
        end else if(((cond_computed5_out & ~cond_stored5_out) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_computed5_write_en = 1'd1;
        end else cond_computed5_write_en = 1'd0;
        cond_computed6_clk = clk;
        if((((~cond_computed6_out & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_in = 1'd1;
        end else if((((cond_stored6_out & cond_computed6_out) & (fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_in = 1'd0;
        end else if(((cond_computed6_out & ~cond_stored6_out) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_in = 1'd0;
        end else cond_computed6_in = 1'd0;
        if((((~cond_computed6_out & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_write_en = 1'd1;
        end else if((((cond_stored6_out & cond_computed6_out) & (fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_write_en = 1'd1;
        end else if(((cond_computed6_out & ~cond_stored6_out) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_write_en = 1'd1;
        end else cond_computed6_write_en = 1'd0;
        cond_computed7_clk = clk;
        if((((~cond_computed7_out & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_in = 1'd1;
        end else if((((cond_stored7_out & cond_computed7_out) & (fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_in = 1'd0;
        end else if(((cond_computed7_out & ~cond_stored7_out) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_in = 1'd0;
        end else cond_computed7_in = 1'd0;
        if((((~cond_computed7_out & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_write_en = 1'd1;
        end else if((((cond_stored7_out & cond_computed7_out) & (fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_write_en = 1'd1;
        end else if(((cond_computed7_out & ~cond_stored7_out) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_write_en = 1'd1;
        end else cond_computed7_write_en = 1'd0;
        cond_computed8_clk = clk;
        if((((~cond_computed8_out & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_in = 1'd1;
        end else if((((cond_stored8_out & cond_computed8_out) & (fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_in = 1'd0;
        end else if(((cond_computed8_out & ~cond_stored8_out) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_in = 1'd0;
        end else cond_computed8_in = 1'd0;
        if((((~cond_computed8_out & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_write_en = 1'd1;
        end else if((((cond_stored8_out & cond_computed8_out) & (fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_write_en = 1'd1;
        end else if(((cond_computed8_out & ~cond_stored8_out) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_write_en = 1'd1;
        end else cond_computed8_write_en = 1'd0;
        cond_computed9_clk = clk;
        if((((~cond_computed9_out & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed9_in = 1'd1;
        end else if((((cond_stored9_out & cond_computed9_out) & (fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed9_in = 1'd0;
        end else if(((cond_computed9_out & ~cond_stored9_out) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed9_in = 1'd0;
        end else cond_computed9_in = 1'd0;
        if((((~cond_computed9_out & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed9_write_en = 1'd1;
        end else if((((cond_stored9_out & cond_computed9_out) & (fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed9_write_en = 1'd1;
        end else if(((cond_computed9_out & ~cond_stored9_out) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_computed9_write_en = 1'd1;
        end else cond_computed9_write_en = 1'd0;
        cond_stored_clk = clk;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_stored_in = le1_out;
        end else cond_stored_in = 1'd0;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_stored_write_en = 1'd1;
        end else cond_stored_write_en = 1'd0;
        cond_stored0_clk = clk;
        if((((~cond_computed0_out & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_stored0_in = le0_out;
        end else cond_stored0_in = 1'd0;
        if((((~cond_computed0_out & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            cond_stored0_write_en = 1'd1;
        end else cond_stored0_write_en = 1'd0;
        cond_stored1_clk = clk;
        if((((~cond_computed1_out & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_stored1_in = le0_out;
        end else cond_stored1_in = 1'd0;
        if((((~cond_computed1_out & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            cond_stored1_write_en = 1'd1;
        end else cond_stored1_write_en = 1'd0;
        cond_stored10_clk = clk;
        if((((~cond_computed10_out & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) & 1'b1) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_stored10_in = le0_out;
        end else cond_stored10_in = 1'd0;
        if((((~cond_computed10_out & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) & 1'b1) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            cond_stored10_write_en = 1'd1;
        end else cond_stored10_write_en = 1'd0;
        cond_stored11_clk = clk;
        if((((~cond_computed11_out & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_stored11_in = le0_out;
        end else cond_stored11_in = 1'd0;
        if((((~cond_computed11_out & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_stored11_write_en = 1'd1;
        end else cond_stored11_write_en = 1'd0;
        cond_stored2_clk = clk;
        if((((~cond_computed2_out & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_stored2_in = le0_out;
        end else cond_stored2_in = 1'd0;
        if((((~cond_computed2_out & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            cond_stored2_write_en = 1'd1;
        end else cond_stored2_write_en = 1'd0;
        cond_stored3_clk = clk;
        if((((~cond_computed3_out & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_stored3_in = le0_out;
        end else cond_stored3_in = 1'd0;
        if((((~cond_computed3_out & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            cond_stored3_write_en = 1'd1;
        end else cond_stored3_write_en = 1'd0;
        cond_stored4_clk = clk;
        if((((~cond_computed4_out & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_stored4_in = le0_out;
        end else cond_stored4_in = 1'd0;
        if((((~cond_computed4_out & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            cond_stored4_write_en = 1'd1;
        end else cond_stored4_write_en = 1'd0;
        cond_stored5_clk = clk;
        if((((~cond_computed5_out & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_stored5_in = le0_out;
        end else cond_stored5_in = 1'd0;
        if((((~cond_computed5_out & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            cond_stored5_write_en = 1'd1;
        end else cond_stored5_write_en = 1'd0;
        cond_stored6_clk = clk;
        if((((~cond_computed6_out & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_stored6_in = le0_out;
        end else cond_stored6_in = 1'd0;
        if((((~cond_computed6_out & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            cond_stored6_write_en = 1'd1;
        end else cond_stored6_write_en = 1'd0;
        cond_stored7_clk = clk;
        if((((~cond_computed7_out & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_stored7_in = le0_out;
        end else cond_stored7_in = 1'd0;
        if((((~cond_computed7_out & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            cond_stored7_write_en = 1'd1;
        end else cond_stored7_write_en = 1'd0;
        cond_stored8_clk = clk;
        if((((~cond_computed8_out & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_stored8_in = le0_out;
        end else cond_stored8_in = 1'd0;
        if((((~cond_computed8_out & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            cond_stored8_write_en = 1'd1;
        end else cond_stored8_write_en = 1'd0;
        cond_stored9_clk = clk;
        if((((~cond_computed9_out & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_stored9_in = le1_out;
        end else cond_stored9_in = 1'd0;
        if((((~cond_computed9_out & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) & 1'b1) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            cond_stored9_write_en = 1'd1;
        end else cond_stored9_write_en = 1'd0;
        done_reg_clk = clk;
        if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            done_reg_in = 1'd1;
        end else if(done_reg_out) begin
            done_reg_in = 1'd0;
        end else done_reg_in = 1'd0;
        if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            done_reg_write_en = 1'd1;
        end else if(done_reg_out) begin
            done_reg_write_en = 1'd1;
        end else done_reg_write_en = 1'd0;
        done_reg0_clk = clk;
        if(((cond_computed0_out & ~cond_stored0_out) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            done_reg0_in = 1'd1;
        end else if(done_reg0_out) begin
            done_reg0_in = 1'd0;
        end else done_reg0_in = 1'd0;
        if(((cond_computed0_out & ~cond_stored0_out) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            done_reg0_write_en = 1'd1;
        end else if(done_reg0_out) begin
            done_reg0_write_en = 1'd1;
        end else done_reg0_write_en = 1'd0;
        done_reg1_clk = clk;
        if(((cond_computed1_out & ~cond_stored1_out) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            done_reg1_in = 1'd1;
        end else if(done_reg1_out) begin
            done_reg1_in = 1'd0;
        end else done_reg1_in = 1'd0;
        if(((cond_computed1_out & ~cond_stored1_out) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            done_reg1_write_en = 1'd1;
        end else if(done_reg1_out) begin
            done_reg1_write_en = 1'd1;
        end else done_reg1_write_en = 1'd0;
        done_reg10_clk = clk;
        if(((cond_computed10_out & ~cond_stored10_out) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            done_reg10_in = 1'd1;
        end else if(done_reg10_out) begin
            done_reg10_in = 1'd0;
        end else done_reg10_in = 1'd0;
        if(((cond_computed10_out & ~cond_stored10_out) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            done_reg10_write_en = 1'd1;
        end else if(done_reg10_out) begin
            done_reg10_write_en = 1'd1;
        end else done_reg10_write_en = 1'd0;
        done_reg11_clk = clk;
        if(((cond_computed11_out & ~cond_stored11_out) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            done_reg11_in = 1'd1;
        end else if(done_reg11_out) begin
            done_reg11_in = 1'd0;
        end else done_reg11_in = 1'd0;
        if(((cond_computed11_out & ~cond_stored11_out) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            done_reg11_write_en = 1'd1;
        end else if(done_reg11_out) begin
            done_reg11_write_en = 1'd1;
        end else done_reg11_write_en = 1'd0;
        done_reg2_clk = clk;
        if(((cond_computed2_out & ~cond_stored2_out) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            done_reg2_in = 1'd1;
        end else if(done_reg2_out) begin
            done_reg2_in = 1'd0;
        end else done_reg2_in = 1'd0;
        if(((cond_computed2_out & ~cond_stored2_out) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            done_reg2_write_en = 1'd1;
        end else if(done_reg2_out) begin
            done_reg2_write_en = 1'd1;
        end else done_reg2_write_en = 1'd0;
        done_reg3_clk = clk;
        if(((cond_computed3_out & ~cond_stored3_out) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            done_reg3_in = 1'd1;
        end else if(done_reg3_out) begin
            done_reg3_in = 1'd0;
        end else done_reg3_in = 1'd0;
        if(((cond_computed3_out & ~cond_stored3_out) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            done_reg3_write_en = 1'd1;
        end else if(done_reg3_out) begin
            done_reg3_write_en = 1'd1;
        end else done_reg3_write_en = 1'd0;
        done_reg4_clk = clk;
        if(((cond_computed4_out & ~cond_stored4_out) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            done_reg4_in = 1'd1;
        end else if(done_reg4_out) begin
            done_reg4_in = 1'd0;
        end else done_reg4_in = 1'd0;
        if(((cond_computed4_out & ~cond_stored4_out) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            done_reg4_write_en = 1'd1;
        end else if(done_reg4_out) begin
            done_reg4_write_en = 1'd1;
        end else done_reg4_write_en = 1'd0;
        done_reg5_clk = clk;
        if(((cond_computed5_out & ~cond_stored5_out) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            done_reg5_in = 1'd1;
        end else if(done_reg5_out) begin
            done_reg5_in = 1'd0;
        end else done_reg5_in = 1'd0;
        if(((cond_computed5_out & ~cond_stored5_out) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            done_reg5_write_en = 1'd1;
        end else if(done_reg5_out) begin
            done_reg5_write_en = 1'd1;
        end else done_reg5_write_en = 1'd0;
        done_reg6_clk = clk;
        if(((cond_computed6_out & ~cond_stored6_out) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            done_reg6_in = 1'd1;
        end else if(done_reg6_out) begin
            done_reg6_in = 1'd0;
        end else done_reg6_in = 1'd0;
        if(((cond_computed6_out & ~cond_stored6_out) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            done_reg6_write_en = 1'd1;
        end else if(done_reg6_out) begin
            done_reg6_write_en = 1'd1;
        end else done_reg6_write_en = 1'd0;
        done_reg7_clk = clk;
        if(((cond_computed7_out & ~cond_stored7_out) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            done_reg7_in = 1'd1;
        end else if(done_reg7_out) begin
            done_reg7_in = 1'd0;
        end else done_reg7_in = 1'd0;
        if(((cond_computed7_out & ~cond_stored7_out) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            done_reg7_write_en = 1'd1;
        end else if(done_reg7_out) begin
            done_reg7_write_en = 1'd1;
        end else done_reg7_write_en = 1'd0;
        done_reg8_clk = clk;
        if(((cond_computed8_out & ~cond_stored8_out) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            done_reg8_in = 1'd1;
        end else if(done_reg8_out) begin
            done_reg8_in = 1'd0;
        end else done_reg8_in = 1'd0;
        if(((cond_computed8_out & ~cond_stored8_out) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            done_reg8_write_en = 1'd1;
        end else if(done_reg8_out) begin
            done_reg8_write_en = 1'd1;
        end else done_reg8_write_en = 1'd0;
        done_reg9_clk = clk;
        if(((cond_computed9_out & ~cond_stored9_out) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            done_reg9_in = 1'd1;
        end else if(done_reg9_out) begin
            done_reg9_in = 1'd0;
        end else done_reg9_in = 1'd0;
        if(((cond_computed9_out & ~cond_stored9_out) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            done_reg9_write_en = 1'd1;
        end else if(done_reg9_out) begin
            done_reg9_write_en = 1'd1;
        end else done_reg9_write_en = 1'd0;
        fsm_clk = clk;
        if((((fsm_out == 32'd0) & u1_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd1;
        end else if((((fsm_out == 32'd1) & par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd2;
        end else if((((fsm_out == 32'd2) & par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd3;
        end else if((((fsm_out == 32'd3) & par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd4;
        end else if((((fsm_out == 32'd4) & par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd5;
        end else if((((fsm_out == 32'd5) & par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd6;
        end else if((((fsm_out == 32'd6) & par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd7;
        end else if((((fsm_out == 32'd7) & par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd8;
        end else if((((fsm_out == 32'd8) & z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd9;
        end else if((((fsm_out == 32'd9) & i0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_in = 32'd10;
        end else if((fsm_out == 32'd10)) begin
            fsm_in = 32'd0;
        end else fsm_in = 32'd0;
        if((((fsm_out == 32'd0) & u1_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd1) & par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd2) & par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd3) & par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd4) & par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd5) & par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd6) & par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd7) & par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd8) & z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd9) & i0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((fsm_out == 32'd10)) begin
            fsm_write_en = 1'd1;
        end else fsm_write_en = 1'd0;
        fsm0_clk = clk;
        if((((fsm0_out == 32'd0) & i0_done) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm0_in = 32'd1;
        end else if((((fsm0_out == 32'd1) & done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm0_in = 32'd2;
        end else if((fsm0_out == 32'd2)) begin
            fsm0_in = 32'd0;
        end else fsm0_in = 32'd0;
        if((((fsm0_out == 32'd0) & i0_done) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm0_write_en = 1'd1;
        end else if((((fsm0_out == 32'd1) & done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm0_write_en = 1'd1;
        end else if((fsm0_out == 32'd2)) begin
            fsm0_write_en = 1'd1;
        end else fsm0_write_en = 1'd0;
        fsm1_clk = clk;
        if((((fsm1_out == 32'd0) & A_int_read0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            fsm1_in = 32'd1;
        end else if((((fsm1_out == 32'd1) & A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            fsm1_in = 32'd2;
        end else if((((fsm1_out == 32'd2) & j0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            fsm1_in = 32'd3;
        end else if((fsm1_out == 32'd3)) begin
            fsm1_in = 32'd0;
        end else fsm1_in = 32'd0;
        if((((fsm1_out == 32'd0) & A_int_read0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd1) & A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd2) & j0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((fsm1_out == 32'd3)) begin
            fsm1_write_en = 1'd1;
        end else fsm1_write_en = 1'd0;
        fsm10_clk = clk;
        if((((fsm10_out == 32'd0) & par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_in = 32'd1;
        end else if((((fsm10_out == 32'd1) & bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_in = 32'd2;
        end else if((((fsm10_out == 32'd2) & bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_in = 32'd3;
        end else if((((fsm10_out == 32'd3) & tmp4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_in = 32'd4;
        end else if((((fsm10_out == 32'd4) & w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_in = 32'd5;
        end else if((((fsm10_out == 32'd5) & j3_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_in = 32'd6;
        end else if((fsm10_out == 32'd6)) begin
            fsm10_in = 32'd0;
        end else fsm10_in = 32'd0;
        if((((fsm10_out == 32'd0) & par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_write_en = 1'd1;
        end else if((((fsm10_out == 32'd1) & bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_write_en = 1'd1;
        end else if((((fsm10_out == 32'd2) & bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_write_en = 1'd1;
        end else if((((fsm10_out == 32'd3) & tmp4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_write_en = 1'd1;
        end else if((((fsm10_out == 32'd4) & w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_write_en = 1'd1;
        end else if((((fsm10_out == 32'd5) & j3_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            fsm10_write_en = 1'd1;
        end else if((fsm10_out == 32'd6)) begin
            fsm10_write_en = 1'd1;
        end else fsm10_write_en = 1'd0;
        fsm11_clk = clk;
        if((((fsm11_out == 32'd0) & j3_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            fsm11_in = 32'd1;
        end else if((((fsm11_out == 32'd1) & done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            fsm11_in = 32'd2;
        end else if((((fsm11_out == 32'd2) & i5_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            fsm11_in = 32'd3;
        end else if((fsm11_out == 32'd3)) begin
            fsm11_in = 32'd0;
        end else fsm11_in = 32'd0;
        if((((fsm11_out == 32'd0) & j3_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            fsm11_write_en = 1'd1;
        end else if((((fsm11_out == 32'd1) & done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            fsm11_write_en = 1'd1;
        end else if((((fsm11_out == 32'd2) & i5_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            fsm11_write_en = 1'd1;
        end else if((fsm11_out == 32'd3)) begin
            fsm11_write_en = 1'd1;
        end else fsm11_write_en = 1'd0;
        fsm12_clk = clk;
        if((((fsm12_out == 32'd0) & u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd1;
        end else if((((fsm12_out == 32'd1) & par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd2;
        end else if((((fsm12_out == 32'd2) & par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd3;
        end else if((((fsm12_out == 32'd3) & par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd4;
        end else if((((fsm12_out == 32'd4) & par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd5;
        end else if((((fsm12_out == 32'd5) & par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd6;
        end else if((((fsm12_out == 32'd6) & par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd7;
        end else if((((fsm12_out == 32'd7) & par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd8;
        end else if((((fsm12_out == 32'd8) & z_int0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd9;
        end else if((((fsm12_out == 32'd9) & i6_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_in = 32'd10;
        end else if((fsm12_out == 32'd10)) begin
            fsm12_in = 32'd0;
        end else fsm12_in = 32'd0;
        if((((fsm12_out == 32'd0) & u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd1) & par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd2) & par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd3) & par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd4) & par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd5) & par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd6) & par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd7) & par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd8) & z_int0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((((fsm12_out == 32'd9) & i6_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm12_write_en = 1'd1;
        end else if((fsm12_out == 32'd10)) begin
            fsm12_write_en = 1'd1;
        end else fsm12_write_en = 1'd0;
        fsm13_clk = clk;
        if((((fsm13_out == 32'd0) & i6_done) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm13_in = 32'd1;
        end else if((((fsm13_out == 32'd1) & done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm13_in = 32'd2;
        end else if((fsm13_out == 32'd2)) begin
            fsm13_in = 32'd0;
        end else fsm13_in = 32'd0;
        if((((fsm13_out == 32'd0) & i6_done) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm13_write_en = 1'd1;
        end else if((((fsm13_out == 32'd1) & done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm13_write_en = 1'd1;
        end else if((fsm13_out == 32'd2)) begin
            fsm13_write_en = 1'd1;
        end else fsm13_write_en = 1'd0;
        fsm14_clk = clk;
        if((((fsm14_out == 32'd0) & A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            fsm14_in = 32'd1;
        end else if((((fsm14_out == 32'd1) & A_int0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            fsm14_in = 32'd2;
        end else if((((fsm14_out == 32'd2) & j4_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            fsm14_in = 32'd3;
        end else if((fsm14_out == 32'd3)) begin
            fsm14_in = 32'd0;
        end else fsm14_in = 32'd0;
        if((((fsm14_out == 32'd0) & A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            fsm14_write_en = 1'd1;
        end else if((((fsm14_out == 32'd1) & A_int0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            fsm14_write_en = 1'd1;
        end else if((((fsm14_out == 32'd2) & j4_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            fsm14_write_en = 1'd1;
        end else if((fsm14_out == 32'd3)) begin
            fsm14_write_en = 1'd1;
        end else fsm14_write_en = 1'd0;
        fsm15_clk = clk;
        if((((fsm15_out == 32'd0) & j4_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm15_in = 32'd1;
        end else if((((fsm15_out == 32'd1) & done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm15_in = 32'd2;
        end else if((((fsm15_out == 32'd2) & i7_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm15_in = 32'd3;
        end else if((fsm15_out == 32'd3)) begin
            fsm15_in = 32'd0;
        end else fsm15_in = 32'd0;
        if((((fsm15_out == 32'd0) & j4_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm15_write_en = 1'd1;
        end else if((((fsm15_out == 32'd1) & done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm15_write_en = 1'd1;
        end else if((((fsm15_out == 32'd2) & i7_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            fsm15_write_en = 1'd1;
        end else if((fsm15_out == 32'd3)) begin
            fsm15_write_en = 1'd1;
        end else fsm15_write_en = 1'd0;
        fsm16_clk = clk;
        if((((fsm16_out == 32'd0) & i7_done) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm16_in = 32'd1;
        end else if((((fsm16_out == 32'd1) & done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm16_in = 32'd2;
        end else if((fsm16_out == 32'd2)) begin
            fsm16_in = 32'd0;
        end else fsm16_in = 32'd0;
        if((((fsm16_out == 32'd0) & i7_done) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm16_write_en = 1'd1;
        end else if((((fsm16_out == 32'd1) & done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            fsm16_write_en = 1'd1;
        end else if((fsm16_out == 32'd2)) begin
            fsm16_write_en = 1'd1;
        end else fsm16_write_en = 1'd0;
        fsm17_clk = clk;
        if((((fsm17_out == 32'd0) & par_reset6_out) & (go | go))) begin
            fsm17_in = 32'd1;
        end else if((((fsm17_out == 32'd1) & i2_done) & (go | go))) begin
            fsm17_in = 32'd2;
        end else if((((fsm17_out == 32'd2) & done_reg3_out) & (go | go))) begin
            fsm17_in = 32'd3;
        end else if((((fsm17_out == 32'd3) & i3_done) & (go | go))) begin
            fsm17_in = 32'd4;
        end else if((((fsm17_out == 32'd4) & done_reg5_out) & (go | go))) begin
            fsm17_in = 32'd5;
        end else if((((fsm17_out == 32'd5) & i4_done) & (go | go))) begin
            fsm17_in = 32'd6;
        end else if((((fsm17_out == 32'd6) & done_reg6_out) & (go | go))) begin
            fsm17_in = 32'd7;
        end else if((((fsm17_out == 32'd7) & i5_done) & (go | go))) begin
            fsm17_in = 32'd8;
        end else if((((fsm17_out == 32'd8) & done_reg8_out) & (go | go))) begin
            fsm17_in = 32'd9;
        end else if((((fsm17_out == 32'd9) & par_reset19_out) & (go | go))) begin
            fsm17_in = 32'd10;
        end else if((fsm17_out == 32'd10)) begin
            fsm17_in = 32'd0;
        end else fsm17_in = 32'd0;
        if((((fsm17_out == 32'd0) & par_reset6_out) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd1) & i2_done) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd2) & done_reg3_out) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd3) & i3_done) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd4) & done_reg5_out) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd5) & i4_done) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd6) & done_reg6_out) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd7) & i5_done) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd8) & done_reg8_out) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((((fsm17_out == 32'd9) & par_reset19_out) & (go | go))) begin
            fsm17_write_en = 1'd1;
        end else if((fsm17_out == 32'd10)) begin
            fsm17_write_en = 1'd1;
        end else fsm17_write_en = 1'd0;
        fsm2_clk = clk;
        if((((fsm2_out == 32'd0) & j0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm2_in = 32'd1;
        end else if((((fsm2_out == 32'd1) & done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm2_in = 32'd2;
        end else if((((fsm2_out == 32'd2) & i1_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm2_in = 32'd3;
        end else if((fsm2_out == 32'd3)) begin
            fsm2_in = 32'd0;
        end else fsm2_in = 32'd0;
        if((((fsm2_out == 32'd0) & j0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((((fsm2_out == 32'd1) & done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((((fsm2_out == 32'd2) & i1_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((fsm2_out == 32'd3)) begin
            fsm2_write_en = 1'd1;
        end else fsm2_write_en = 1'd0;
        fsm3_clk = clk;
        if((((fsm3_out == 32'd0) & i1_done) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm3_in = 32'd1;
        end else if((((fsm3_out == 32'd1) & done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm3_in = 32'd2;
        end else if((fsm3_out == 32'd2)) begin
            fsm3_in = 32'd0;
        end else fsm3_in = 32'd0;
        if((((fsm3_out == 32'd0) & i1_done) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm3_write_en = 1'd1;
        end else if((((fsm3_out == 32'd1) & done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            fsm3_write_en = 1'd1;
        end else if((fsm3_out == 32'd2)) begin
            fsm3_write_en = 1'd1;
        end else fsm3_write_en = 1'd0;
        fsm4_clk = clk;
        if((((fsm4_out == 32'd0) & bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            fsm4_in = 32'd1;
        end else if((((fsm4_out == 32'd1) & bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            fsm4_in = 32'd2;
        end else if((((fsm4_out == 32'd2) & tmp1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            fsm4_in = 32'd3;
        end else if((fsm4_out == 32'd3)) begin
            fsm4_in = 32'd0;
        end else fsm4_in = 32'd0;
        if((((fsm4_out == 32'd0) & bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((((fsm4_out == 32'd1) & bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((((fsm4_out == 32'd2) & tmp1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((fsm4_out == 32'd3)) begin
            fsm4_write_en = 1'd1;
        end else fsm4_write_en = 1'd0;
        fsm5_clk = clk;
        if((((fsm5_out == 32'd0) & par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_in = 32'd1;
        end else if((((fsm5_out == 32'd1) & par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_in = 32'd2;
        end else if((((fsm5_out == 32'd2) & A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_in = 32'd3;
        end else if((((fsm5_out == 32'd3) & j1_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_in = 32'd4;
        end else if((fsm5_out == 32'd4)) begin
            fsm5_in = 32'd0;
        end else fsm5_in = 32'd0;
        if((((fsm5_out == 32'd0) & par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd1) & par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd2) & A0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd3) & j1_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((fsm5_out == 32'd4)) begin
            fsm5_write_en = 1'd1;
        end else fsm5_write_en = 1'd0;
        fsm6_clk = clk;
        if((((fsm6_out == 32'd0) & j1_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            fsm6_in = 32'd1;
        end else if((((fsm6_out == 32'd1) & done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            fsm6_in = 32'd2;
        end else if((((fsm6_out == 32'd2) & i2_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            fsm6_in = 32'd3;
        end else if((fsm6_out == 32'd3)) begin
            fsm6_in = 32'd0;
        end else fsm6_in = 32'd0;
        if((((fsm6_out == 32'd0) & j1_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            fsm6_write_en = 1'd1;
        end else if((((fsm6_out == 32'd1) & done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            fsm6_write_en = 1'd1;
        end else if((((fsm6_out == 32'd2) & i2_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            fsm6_write_en = 1'd1;
        end else if((fsm6_out == 32'd3)) begin
            fsm6_write_en = 1'd1;
        end else fsm6_write_en = 1'd0;
        fsm7_clk = clk;
        if((((fsm7_out == 32'd0) & par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_in = 32'd1;
        end else if((((fsm7_out == 32'd1) & bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_in = 32'd2;
        end else if((((fsm7_out == 32'd2) & bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_in = 32'd3;
        end else if((((fsm7_out == 32'd3) & tmp2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_in = 32'd4;
        end else if((((fsm7_out == 32'd4) & x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_in = 32'd5;
        end else if((((fsm7_out == 32'd5) & j2_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_in = 32'd6;
        end else if((fsm7_out == 32'd6)) begin
            fsm7_in = 32'd0;
        end else fsm7_in = 32'd0;
        if((((fsm7_out == 32'd0) & par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd1) & bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd2) & bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd3) & tmp2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd4) & x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd5) & j2_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((fsm7_out == 32'd6)) begin
            fsm7_write_en = 1'd1;
        end else fsm7_write_en = 1'd0;
        fsm8_clk = clk;
        if((((fsm8_out == 32'd0) & j2_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            fsm8_in = 32'd1;
        end else if((((fsm8_out == 32'd1) & done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            fsm8_in = 32'd2;
        end else if((((fsm8_out == 32'd2) & i3_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            fsm8_in = 32'd3;
        end else if((fsm8_out == 32'd3)) begin
            fsm8_in = 32'd0;
        end else fsm8_in = 32'd0;
        if((((fsm8_out == 32'd0) & j2_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            fsm8_write_en = 1'd1;
        end else if((((fsm8_out == 32'd1) & done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            fsm8_write_en = 1'd1;
        end else if((((fsm8_out == 32'd2) & i3_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            fsm8_write_en = 1'd1;
        end else if((fsm8_out == 32'd3)) begin
            fsm8_write_en = 1'd1;
        end else fsm8_write_en = 1'd0;
        fsm9_clk = clk;
        if((((fsm9_out == 32'd0) & par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            fsm9_in = 32'd1;
        end else if((((fsm9_out == 32'd1) & x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            fsm9_in = 32'd2;
        end else if((((fsm9_out == 32'd2) & i4_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            fsm9_in = 32'd3;
        end else if((fsm9_out == 32'd3)) begin
            fsm9_in = 32'd0;
        end else fsm9_in = 32'd0;
        if((((fsm9_out == 32'd0) & par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd1) & x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd2) & i4_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            fsm9_write_en = 1'd1;
        end else if((fsm9_out == 32'd3)) begin
            fsm9_write_en = 1'd1;
        end else fsm9_write_en = 1'd0;
        i0_clk = clk;
        if((((fsm0_out == 32'd0) & ~i0_done) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            i0_in = const13_out;
        end else if((((fsm_out == 32'd9) & ~i0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            i0_in = add1_out;
        end else i0_in = 7'd0;
        if((((fsm0_out == 32'd0) & ~i0_done) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            i0_write_en = 1'd1;
        end else if((((fsm_out == 32'd9) & ~i0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            i0_write_en = 1'd1;
        end else i0_write_en = 1'd0;
        i1_clk = clk;
        if((((fsm3_out == 32'd0) & ~i1_done) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            i1_in = const10_out;
        end else if((((fsm2_out == 32'd2) & ~i1_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            i1_in = add0_out;
        end else i1_in = 7'd0;
        if((((fsm3_out == 32'd0) & ~i1_done) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))) begin
            i1_write_en = 1'd1;
        end else if((((fsm2_out == 32'd2) & ~i1_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            i1_write_en = 1'd1;
        end else i1_write_en = 1'd0;
        i2_clk = clk;
        if((((fsm17_out == 32'd1) & ~i2_done) & (go | go))) begin
            i2_in = const10_out;
        end else if((((fsm6_out == 32'd2) & ~i2_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            i2_in = add0_out;
        end else i2_in = 7'd0;
        if((((fsm17_out == 32'd1) & ~i2_done) & (go | go))) begin
            i2_write_en = 1'd1;
        end else if((((fsm6_out == 32'd2) & ~i2_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            i2_write_en = 1'd1;
        end else i2_write_en = 1'd0;
        i3_clk = clk;
        if((((fsm17_out == 32'd3) & ~i3_done) & (go | go))) begin
            i3_in = const10_out;
        end else if((((fsm8_out == 32'd2) & ~i3_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            i3_in = add0_out;
        end else i3_in = 7'd0;
        if((((fsm17_out == 32'd3) & ~i3_done) & (go | go))) begin
            i3_write_en = 1'd1;
        end else if((((fsm8_out == 32'd2) & ~i3_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            i3_write_en = 1'd1;
        end else i3_write_en = 1'd0;
        i4_clk = clk;
        if((((fsm17_out == 32'd5) & ~i4_done) & (go | go))) begin
            i4_in = const10_out;
        end else if((((fsm9_out == 32'd2) & ~i4_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            i4_in = add0_out;
        end else i4_in = 7'd0;
        if((((fsm17_out == 32'd5) & ~i4_done) & (go | go))) begin
            i4_write_en = 1'd1;
        end else if((((fsm9_out == 32'd2) & ~i4_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            i4_write_en = 1'd1;
        end else i4_write_en = 1'd0;
        i5_clk = clk;
        if((((fsm17_out == 32'd7) & ~i5_done) & (go | go))) begin
            i5_in = const10_out;
        end else if((((fsm11_out == 32'd2) & ~i5_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            i5_in = add0_out;
        end else i5_in = 7'd0;
        if((((fsm17_out == 32'd7) & ~i5_done) & (go | go))) begin
            i5_write_en = 1'd1;
        end else if((((fsm11_out == 32'd2) & ~i5_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            i5_write_en = 1'd1;
        end else i5_write_en = 1'd0;
        i6_clk = clk;
        if((((fsm13_out == 32'd0) & ~i6_done) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            i6_in = const13_out;
        end else if((((fsm12_out == 32'd9) & ~i6_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            i6_in = add1_out;
        end else i6_in = 7'd0;
        if((((fsm13_out == 32'd0) & ~i6_done) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            i6_write_en = 1'd1;
        end else if((((fsm12_out == 32'd9) & ~i6_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            i6_write_en = 1'd1;
        end else i6_write_en = 1'd0;
        i7_clk = clk;
        if((((fsm16_out == 32'd0) & ~i7_done) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            i7_in = const10_out;
        end else if((((fsm15_out == 32'd2) & ~i7_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            i7_in = add0_out;
        end else i7_in = 7'd0;
        if((((fsm16_out == 32'd0) & ~i7_done) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))) begin
            i7_write_en = 1'd1;
        end else if((((fsm15_out == 32'd2) & ~i7_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            i7_write_en = 1'd1;
        end else i7_write_en = 1'd0;
        j0_clk = clk;
        if((((fsm2_out == 32'd0) & ~j0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            j0_in = const10_out;
        end else if((((fsm1_out == 32'd2) & ~j0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            j0_in = add0_out;
        end else j0_in = 7'd0;
        if((((fsm2_out == 32'd0) & ~j0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            j0_write_en = 1'd1;
        end else if((((fsm1_out == 32'd2) & ~j0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            j0_write_en = 1'd1;
        end else j0_write_en = 1'd0;
        j1_clk = clk;
        if((((fsm6_out == 32'd0) & ~j1_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            j1_in = const10_out;
        end else if((((fsm5_out == 32'd3) & ~j1_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            j1_in = add0_out;
        end else j1_in = 7'd0;
        if((((fsm6_out == 32'd0) & ~j1_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))) begin
            j1_write_en = 1'd1;
        end else if((((fsm5_out == 32'd3) & ~j1_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))) begin
            j1_write_en = 1'd1;
        end else j1_write_en = 1'd0;
        j2_clk = clk;
        if((((fsm8_out == 32'd0) & ~j2_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            j2_in = const10_out;
        end else if((((fsm7_out == 32'd5) & ~j2_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            j2_in = add0_out;
        end else j2_in = 7'd0;
        if((((fsm8_out == 32'd0) & ~j2_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))) begin
            j2_write_en = 1'd1;
        end else if((((fsm7_out == 32'd5) & ~j2_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            j2_write_en = 1'd1;
        end else j2_write_en = 1'd0;
        j3_clk = clk;
        if((((fsm11_out == 32'd0) & ~j3_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            j3_in = const10_out;
        end else if((((fsm10_out == 32'd5) & ~j3_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            j3_in = add0_out;
        end else j3_in = 7'd0;
        if((((fsm11_out == 32'd0) & ~j3_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))) begin
            j3_write_en = 1'd1;
        end else if((((fsm10_out == 32'd5) & ~j3_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            j3_write_en = 1'd1;
        end else j3_write_en = 1'd0;
        j4_clk = clk;
        if((((fsm15_out == 32'd0) & ~j4_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            j4_in = const10_out;
        end else if((((fsm14_out == 32'd2) & ~j4_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            j4_in = add0_out;
        end else j4_in = 7'd0;
        if((((fsm15_out == 32'd0) & ~j4_done) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            j4_write_en = 1'd1;
        end else if((((fsm14_out == 32'd2) & ~j4_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            j4_write_en = 1'd1;
        end else j4_write_en = 1'd0;
        if((~cond_computed1_out & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            le0_left = i1_out;
        end else if((~cond_computed11_out & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            le0_left = i7_out;
        end else if((~cond_computed10_out & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            le0_left = j4_out;
        end else if((~cond_computed0_out & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            le0_left = j0_out;
        end else if((~cond_computed3_out & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            le0_left = i2_out;
        end else if((~cond_computed2_out & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            le0_left = j1_out;
        end else if((~cond_computed5_out & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            le0_left = i3_out;
        end else if((~cond_computed4_out & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            le0_left = j2_out;
        end else if((~cond_computed6_out & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            le0_left = i4_out;
        end else if((~cond_computed8_out & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            le0_left = i5_out;
        end else if((~cond_computed7_out & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            le0_left = j3_out;
        end else le0_left = 7'd0;
        if((~cond_computed1_out & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            le0_right = const14_out;
        end else if((~cond_computed11_out & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            le0_right = const14_out;
        end else if((~cond_computed10_out & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            le0_right = const14_out;
        end else if((~cond_computed0_out & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            le0_right = const14_out;
        end else if((~cond_computed3_out & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))) begin
            le0_right = const14_out;
        end else if((~cond_computed2_out & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))) begin
            le0_right = const14_out;
        end else if((~cond_computed5_out & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))) begin
            le0_right = const14_out;
        end else if((~cond_computed4_out & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))) begin
            le0_right = const14_out;
        end else if((~cond_computed6_out & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))) begin
            le0_right = const14_out;
        end else if((~cond_computed8_out & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))) begin
            le0_right = const14_out;
        end else if((~cond_computed7_out & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))) begin
            le0_right = const14_out;
        end else le0_right = 7'd0;
        if((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            le1_left = i0_out;
        end else if((~cond_computed9_out & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            le1_left = i6_out;
        end else le1_left = 7'd0;
        if((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))) begin
            le1_right = const16_out;
        end else if((~cond_computed9_out & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))) begin
            le1_right = const16_out;
        end else le1_right = 7'd0;
        mult_pipe0_clk = clk;
        if((~mult_pipe0_done & (((fsm4_out == 32'd0) & ~bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))))) begin
            mult_pipe0_go = 1'd1;
        end else mult_pipe0_go = 1'd0;
        if((((fsm4_out == 32'd0) & ~bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe0_left = u1_read0_0_out;
        end else mult_pipe0_left = 32'd0;
        if((((fsm4_out == 32'd0) & ~bin_read0_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe0_right = v1_read0_0_out;
        end else mult_pipe0_right = 32'd0;
        mult_pipe1_clk = clk;
        if((~mult_pipe1_done & (((fsm4_out == 32'd1) & ~bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))))) begin
            mult_pipe1_go = 1'd1;
        end else mult_pipe1_go = 1'd0;
        if((((fsm4_out == 32'd1) & ~bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe1_left = u2_read0_0_out;
        end else mult_pipe1_left = 32'd0;
        if((((fsm4_out == 32'd1) & ~bin_read1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe1_right = v2_read0_0_out;
        end else mult_pipe1_right = 32'd0;
        mult_pipe2_clk = clk;
        if((~mult_pipe2_done & (((fsm7_out == 32'd1) & ~bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            mult_pipe2_go = 1'd1;
        end else mult_pipe2_go = 1'd0;
        if((((fsm7_out == 32'd1) & ~bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            mult_pipe2_left = beta__0_out;
        end else mult_pipe2_left = 32'd0;
        if((((fsm7_out == 32'd1) & ~bin_read2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            mult_pipe2_right = A_read0_0_out;
        end else mult_pipe2_right = 32'd0;
        mult_pipe3_clk = clk;
        if((~mult_pipe3_done & (((fsm7_out == 32'd2) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            mult_pipe3_go = 1'd1;
        end else mult_pipe3_go = 1'd0;
        if((((fsm7_out == 32'd2) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            mult_pipe3_left = bin_read2_0_out;
        end else mult_pipe3_left = 32'd0;
        if((((fsm7_out == 32'd2) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            mult_pipe3_right = y_read0_0_out;
        end else mult_pipe3_right = 32'd0;
        mult_pipe4_clk = clk;
        if((~mult_pipe4_done & (((fsm10_out == 32'd1) & ~bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            mult_pipe4_go = 1'd1;
        end else mult_pipe4_go = 1'd0;
        if((((fsm10_out == 32'd1) & ~bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            mult_pipe4_left = alpha__0_out;
        end else mult_pipe4_left = 32'd0;
        if((((fsm10_out == 32'd1) & ~bin_read4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            mult_pipe4_right = A_read1_0_out;
        end else mult_pipe4_right = 32'd0;
        mult_pipe5_clk = clk;
        if((~mult_pipe5_done & (((fsm10_out == 32'd2) & ~bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            mult_pipe5_go = 1'd1;
        end else mult_pipe5_go = 1'd0;
        if((((fsm10_out == 32'd2) & ~bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            mult_pipe5_left = bin_read4_0_out;
        end else mult_pipe5_left = 32'd0;
        if((((fsm10_out == 32'd2) & ~bin_read5_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            mult_pipe5_right = x_read0_0_out;
        end else mult_pipe5_right = 32'd0;
        old_0_clk = clk;
        if((~(par_done_reg22_out | old_0_done) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            old_0_in = A0_0_read_data;
        end else old_0_in = 32'd0;
        if((~(par_done_reg22_out | old_0_done) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            old_0_write_en = 1'd1;
        end else old_0_write_en = 1'd0;
        old_1_clk = clk;
        if((~(par_done_reg26_out | old_1_done) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            old_1_in = x0_read_data;
        end else old_1_in = 32'd0;
        if((~(par_done_reg26_out | old_1_done) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            old_1_write_en = 1'd1;
        end else old_1_write_en = 1'd0;
        par_done_reg_clk = clk;
        if((u10_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg_in = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg_in = 1'd0;
        end else par_done_reg_in = 1'd0;
        if((u10_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg_write_en = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg_write_en = 1'd1;
        end else par_done_reg_write_en = 1'd0;
        par_done_reg0_clk = clk;
        if((v1_int_read0_0_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg0_in = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg0_in = 1'd0;
        end else par_done_reg0_in = 1'd0;
        if((v1_int_read0_0_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg0_write_en = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg0_write_en = 1'd1;
        end else par_done_reg0_write_en = 1'd0;
        par_done_reg1_clk = clk;
        if((v10_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg1_in = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg1_in = 1'd0;
        end else par_done_reg1_in = 1'd0;
        if((v10_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg1_write_en = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg1_write_en = 1'd1;
        end else par_done_reg1_write_en = 1'd0;
        par_done_reg10_clk = clk;
        if((y_int_read0_0_done & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg10_in = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg10_in = 1'd0;
        end else par_done_reg10_in = 1'd0;
        if((y_int_read0_0_done & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg10_write_en = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg10_write_en = 1'd1;
        end else par_done_reg10_write_en = 1'd0;
        par_done_reg11_clk = clk;
        if((y0_done & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg11_in = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg11_in = 1'd0;
        end else par_done_reg11_in = 1'd0;
        if((y0_done & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg11_write_en = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg11_write_en = 1'd1;
        end else par_done_reg11_write_en = 1'd0;
        par_done_reg12_clk = clk;
        if((z_int_read0_0_done & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg12_in = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg12_in = 1'd0;
        end else par_done_reg12_in = 1'd0;
        if((z_int_read0_0_done & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg12_write_en = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg12_write_en = 1'd1;
        end else par_done_reg12_write_en = 1'd0;
        par_done_reg13_clk = clk;
        if((alpha__0_done & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg13_in = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg13_in = 1'd0;
        end else par_done_reg13_in = 1'd0;
        if((alpha__0_done & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg13_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg13_write_en = 1'd1;
        end else par_done_reg13_write_en = 1'd0;
        par_done_reg14_clk = clk;
        if((beta__0_done & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg14_in = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg14_in = 1'd0;
        end else par_done_reg14_in = 1'd0;
        if((beta__0_done & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg14_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg14_write_en = 1'd1;
        end else par_done_reg14_write_en = 1'd0;
        par_done_reg15_clk = clk;
        if(((fsm0_out == 32'd2) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg15_in = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg15_in = 1'd0;
        end else par_done_reg15_in = 1'd0;
        if(((fsm0_out == 32'd2) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg15_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg15_write_en = 1'd1;
        end else par_done_reg15_write_en = 1'd0;
        par_done_reg16_clk = clk;
        if(((fsm3_out == 32'd2) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg16_in = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg16_in = 1'd0;
        end else par_done_reg16_in = 1'd0;
        if(((fsm3_out == 32'd2) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_done_reg16_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg16_write_en = 1'd1;
        end else par_done_reg16_write_en = 1'd0;
        par_done_reg17_clk = clk;
        if((u1_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg17_in = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg17_in = 1'd0;
        end else par_done_reg17_in = 1'd0;
        if((u1_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg17_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg17_write_en = 1'd1;
        end else par_done_reg17_write_en = 1'd0;
        par_done_reg18_clk = clk;
        if((v1_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg18_in = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg18_in = 1'd0;
        end else par_done_reg18_in = 1'd0;
        if((v1_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg18_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg18_write_en = 1'd1;
        end else par_done_reg18_write_en = 1'd0;
        par_done_reg19_clk = clk;
        if((u2_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg19_in = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg19_in = 1'd0;
        end else par_done_reg19_in = 1'd0;
        if((u2_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg19_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg19_write_en = 1'd1;
        end else par_done_reg19_write_en = 1'd0;
        par_done_reg2_clk = clk;
        if((u2_int_read0_0_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg2_in = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg2_in = 1'd0;
        end else par_done_reg2_in = 1'd0;
        if((u2_int_read0_0_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg2_write_en = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg2_write_en = 1'd1;
        end else par_done_reg2_write_en = 1'd0;
        par_done_reg20_clk = clk;
        if((v2_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg20_in = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg20_in = 1'd0;
        end else par_done_reg20_in = 1'd0;
        if((v2_read0_0_done & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg20_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg20_write_en = 1'd1;
        end else par_done_reg20_write_en = 1'd0;
        par_done_reg21_clk = clk;
        if(((fsm4_out == 32'd3) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg21_in = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg21_in = 1'd0;
        end else par_done_reg21_in = 1'd0;
        if(((fsm4_out == 32'd3) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg21_write_en = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg21_write_en = 1'd1;
        end else par_done_reg21_write_en = 1'd0;
        par_done_reg22_clk = clk;
        if((old_0_done & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg22_in = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg22_in = 1'd0;
        end else par_done_reg22_in = 1'd0;
        if((old_0_done & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_done_reg22_write_en = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg22_write_en = 1'd1;
        end else par_done_reg22_write_en = 1'd0;
        par_done_reg23_clk = clk;
        if((A_read0_0_done & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            par_done_reg23_in = 1'd1;
        end else if(par_reset9_out) begin
            par_done_reg23_in = 1'd0;
        end else par_done_reg23_in = 1'd0;
        if((A_read0_0_done & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            par_done_reg23_write_en = 1'd1;
        end else if(par_reset9_out) begin
            par_done_reg23_write_en = 1'd1;
        end else par_done_reg23_write_en = 1'd0;
        par_done_reg24_clk = clk;
        if((y_read0_0_done & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            par_done_reg24_in = 1'd1;
        end else if(par_reset9_out) begin
            par_done_reg24_in = 1'd0;
        end else par_done_reg24_in = 1'd0;
        if((y_read0_0_done & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            par_done_reg24_write_en = 1'd1;
        end else if(par_reset9_out) begin
            par_done_reg24_write_en = 1'd1;
        end else par_done_reg24_write_en = 1'd0;
        par_done_reg25_clk = clk;
        if((tmp3_0_done & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            par_done_reg25_in = 1'd1;
        end else if(par_reset10_out) begin
            par_done_reg25_in = 1'd0;
        end else par_done_reg25_in = 1'd0;
        if((tmp3_0_done & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            par_done_reg25_write_en = 1'd1;
        end else if(par_reset10_out) begin
            par_done_reg25_write_en = 1'd1;
        end else par_done_reg25_write_en = 1'd0;
        par_done_reg26_clk = clk;
        if((old_1_done & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            par_done_reg26_in = 1'd1;
        end else if(par_reset10_out) begin
            par_done_reg26_in = 1'd0;
        end else par_done_reg26_in = 1'd0;
        if((old_1_done & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            par_done_reg26_write_en = 1'd1;
        end else if(par_reset10_out) begin
            par_done_reg26_write_en = 1'd1;
        end else par_done_reg26_write_en = 1'd0;
        par_done_reg27_clk = clk;
        if((A_read1_0_done & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg27_in = 1'd1;
        end else if(par_reset11_out) begin
            par_done_reg27_in = 1'd0;
        end else par_done_reg27_in = 1'd0;
        if((A_read1_0_done & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg27_write_en = 1'd1;
        end else if(par_reset11_out) begin
            par_done_reg27_write_en = 1'd1;
        end else par_done_reg27_write_en = 1'd0;
        par_done_reg28_clk = clk;
        if((x_read0_0_done & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg28_in = 1'd1;
        end else if(par_reset11_out) begin
            par_done_reg28_in = 1'd0;
        end else par_done_reg28_in = 1'd0;
        if((x_read0_0_done & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg28_write_en = 1'd1;
        end else if(par_reset11_out) begin
            par_done_reg28_write_en = 1'd1;
        end else par_done_reg28_write_en = 1'd0;
        par_done_reg29_clk = clk;
        if((u1_int0_done & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg29_in = 1'd1;
        end else if(par_reset12_out) begin
            par_done_reg29_in = 1'd0;
        end else par_done_reg29_in = 1'd0;
        if((u1_int0_done & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg29_write_en = 1'd1;
        end else if(par_reset12_out) begin
            par_done_reg29_write_en = 1'd1;
        end else par_done_reg29_write_en = 1'd0;
        par_done_reg3_clk = clk;
        if((u20_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg3_in = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg3_in = 1'd0;
        end else par_done_reg3_in = 1'd0;
        if((u20_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg3_write_en = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg3_write_en = 1'd1;
        end else par_done_reg3_write_en = 1'd0;
        par_done_reg30_clk = clk;
        if((v1_sh_read0_0_done & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg30_in = 1'd1;
        end else if(par_reset12_out) begin
            par_done_reg30_in = 1'd0;
        end else par_done_reg30_in = 1'd0;
        if((v1_sh_read0_0_done & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg30_write_en = 1'd1;
        end else if(par_reset12_out) begin
            par_done_reg30_write_en = 1'd1;
        end else par_done_reg30_write_en = 1'd0;
        par_done_reg31_clk = clk;
        if((v1_int0_done & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg31_in = 1'd1;
        end else if(par_reset13_out) begin
            par_done_reg31_in = 1'd0;
        end else par_done_reg31_in = 1'd0;
        if((v1_int0_done & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg31_write_en = 1'd1;
        end else if(par_reset13_out) begin
            par_done_reg31_write_en = 1'd1;
        end else par_done_reg31_write_en = 1'd0;
        par_done_reg32_clk = clk;
        if((u2_sh_read0_0_done & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg32_in = 1'd1;
        end else if(par_reset13_out) begin
            par_done_reg32_in = 1'd0;
        end else par_done_reg32_in = 1'd0;
        if((u2_sh_read0_0_done & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg32_write_en = 1'd1;
        end else if(par_reset13_out) begin
            par_done_reg32_write_en = 1'd1;
        end else par_done_reg32_write_en = 1'd0;
        par_done_reg33_clk = clk;
        if((u2_int0_done & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg33_in = 1'd1;
        end else if(par_reset14_out) begin
            par_done_reg33_in = 1'd0;
        end else par_done_reg33_in = 1'd0;
        if((u2_int0_done & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg33_write_en = 1'd1;
        end else if(par_reset14_out) begin
            par_done_reg33_write_en = 1'd1;
        end else par_done_reg33_write_en = 1'd0;
        par_done_reg34_clk = clk;
        if((v2_sh_read0_0_done & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg34_in = 1'd1;
        end else if(par_reset14_out) begin
            par_done_reg34_in = 1'd0;
        end else par_done_reg34_in = 1'd0;
        if((v2_sh_read0_0_done & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg34_write_en = 1'd1;
        end else if(par_reset14_out) begin
            par_done_reg34_write_en = 1'd1;
        end else par_done_reg34_write_en = 1'd0;
        par_done_reg35_clk = clk;
        if((v2_int0_done & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg35_in = 1'd1;
        end else if(par_reset15_out) begin
            par_done_reg35_in = 1'd0;
        end else par_done_reg35_in = 1'd0;
        if((v2_int0_done & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg35_write_en = 1'd1;
        end else if(par_reset15_out) begin
            par_done_reg35_write_en = 1'd1;
        end else par_done_reg35_write_en = 1'd0;
        par_done_reg36_clk = clk;
        if((w_sh_read0_0_done & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg36_in = 1'd1;
        end else if(par_reset15_out) begin
            par_done_reg36_in = 1'd0;
        end else par_done_reg36_in = 1'd0;
        if((w_sh_read0_0_done & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg36_write_en = 1'd1;
        end else if(par_reset15_out) begin
            par_done_reg36_write_en = 1'd1;
        end else par_done_reg36_write_en = 1'd0;
        par_done_reg37_clk = clk;
        if((w_int0_done & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg37_in = 1'd1;
        end else if(par_reset16_out) begin
            par_done_reg37_in = 1'd0;
        end else par_done_reg37_in = 1'd0;
        if((w_int0_done & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg37_write_en = 1'd1;
        end else if(par_reset16_out) begin
            par_done_reg37_write_en = 1'd1;
        end else par_done_reg37_write_en = 1'd0;
        par_done_reg38_clk = clk;
        if((x_sh_read0_0_done & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg38_in = 1'd1;
        end else if(par_reset16_out) begin
            par_done_reg38_in = 1'd0;
        end else par_done_reg38_in = 1'd0;
        if((x_sh_read0_0_done & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg38_write_en = 1'd1;
        end else if(par_reset16_out) begin
            par_done_reg38_write_en = 1'd1;
        end else par_done_reg38_write_en = 1'd0;
        par_done_reg39_clk = clk;
        if((x_int0_done & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg39_in = 1'd1;
        end else if(par_reset17_out) begin
            par_done_reg39_in = 1'd0;
        end else par_done_reg39_in = 1'd0;
        if((x_int0_done & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg39_write_en = 1'd1;
        end else if(par_reset17_out) begin
            par_done_reg39_write_en = 1'd1;
        end else par_done_reg39_write_en = 1'd0;
        par_done_reg4_clk = clk;
        if((v2_int_read0_0_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg4_in = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg4_in = 1'd0;
        end else par_done_reg4_in = 1'd0;
        if((v2_int_read0_0_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg4_write_en = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg4_write_en = 1'd1;
        end else par_done_reg4_write_en = 1'd0;
        par_done_reg40_clk = clk;
        if((y_sh_read0_0_done & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg40_in = 1'd1;
        end else if(par_reset17_out) begin
            par_done_reg40_in = 1'd0;
        end else par_done_reg40_in = 1'd0;
        if((y_sh_read0_0_done & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg40_write_en = 1'd1;
        end else if(par_reset17_out) begin
            par_done_reg40_write_en = 1'd1;
        end else par_done_reg40_write_en = 1'd0;
        par_done_reg41_clk = clk;
        if((y_int0_done & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg41_in = 1'd1;
        end else if(par_reset18_out) begin
            par_done_reg41_in = 1'd0;
        end else par_done_reg41_in = 1'd0;
        if((y_int0_done & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg41_write_en = 1'd1;
        end else if(par_reset18_out) begin
            par_done_reg41_write_en = 1'd1;
        end else par_done_reg41_write_en = 1'd0;
        par_done_reg42_clk = clk;
        if((z_sh_read0_0_done & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg42_in = 1'd1;
        end else if(par_reset18_out) begin
            par_done_reg42_in = 1'd0;
        end else par_done_reg42_in = 1'd0;
        if((z_sh_read0_0_done & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_done_reg42_write_en = 1'd1;
        end else if(par_reset18_out) begin
            par_done_reg42_write_en = 1'd1;
        end else par_done_reg42_write_en = 1'd0;
        par_done_reg43_clk = clk;
        if(((fsm13_out == 32'd2) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))) begin
            par_done_reg43_in = 1'd1;
        end else if(par_reset19_out) begin
            par_done_reg43_in = 1'd0;
        end else par_done_reg43_in = 1'd0;
        if(((fsm13_out == 32'd2) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))) begin
            par_done_reg43_write_en = 1'd1;
        end else if(par_reset19_out) begin
            par_done_reg43_write_en = 1'd1;
        end else par_done_reg43_write_en = 1'd0;
        par_done_reg44_clk = clk;
        if(((fsm16_out == 32'd2) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))) begin
            par_done_reg44_in = 1'd1;
        end else if(par_reset19_out) begin
            par_done_reg44_in = 1'd0;
        end else par_done_reg44_in = 1'd0;
        if(((fsm16_out == 32'd2) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))) begin
            par_done_reg44_write_en = 1'd1;
        end else if(par_reset19_out) begin
            par_done_reg44_write_en = 1'd1;
        end else par_done_reg44_write_en = 1'd0;
        par_done_reg5_clk = clk;
        if((v20_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg5_in = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg5_in = 1'd0;
        end else par_done_reg5_in = 1'd0;
        if((v20_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg5_write_en = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg5_write_en = 1'd1;
        end else par_done_reg5_write_en = 1'd0;
        par_done_reg6_clk = clk;
        if((w_int_read0_0_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg6_in = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg6_in = 1'd0;
        end else par_done_reg6_in = 1'd0;
        if((w_int_read0_0_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg6_write_en = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg6_write_en = 1'd1;
        end else par_done_reg6_write_en = 1'd0;
        par_done_reg7_clk = clk;
        if((w0_done & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg7_in = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg7_in = 1'd0;
        end else par_done_reg7_in = 1'd0;
        if((w0_done & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg7_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg7_write_en = 1'd1;
        end else par_done_reg7_write_en = 1'd0;
        par_done_reg8_clk = clk;
        if((x_int_read0_0_done & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg8_in = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg8_in = 1'd0;
        end else par_done_reg8_in = 1'd0;
        if((x_int_read0_0_done & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg8_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg8_write_en = 1'd1;
        end else par_done_reg8_write_en = 1'd0;
        par_done_reg9_clk = clk;
        if((x0_done & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg9_in = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg9_in = 1'd0;
        end else par_done_reg9_in = 1'd0;
        if((x0_done & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_done_reg9_write_en = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg9_write_en = 1'd1;
        end else par_done_reg9_write_en = 1'd0;
        par_reset_clk = clk;
        if(((par_done_reg_out & par_done_reg0_out) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset_in = 1'd1;
        end else if(par_reset_out) begin
            par_reset_in = 1'd0;
        end else par_reset_in = 1'd0;
        if(((par_done_reg_out & par_done_reg0_out) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset_write_en = 1'd1;
        end else if(par_reset_out) begin
            par_reset_write_en = 1'd1;
        end else par_reset_write_en = 1'd0;
        par_reset0_clk = clk;
        if(((par_done_reg1_out & par_done_reg2_out) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset0_in = 1'd1;
        end else if(par_reset0_out) begin
            par_reset0_in = 1'd0;
        end else par_reset0_in = 1'd0;
        if(((par_done_reg1_out & par_done_reg2_out) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset0_write_en = 1'd1;
        end else if(par_reset0_out) begin
            par_reset0_write_en = 1'd1;
        end else par_reset0_write_en = 1'd0;
        par_reset1_clk = clk;
        if(((par_done_reg3_out & par_done_reg4_out) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset1_in = 1'd1;
        end else if(par_reset1_out) begin
            par_reset1_in = 1'd0;
        end else par_reset1_in = 1'd0;
        if(((par_done_reg3_out & par_done_reg4_out) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset1_write_en = 1'd1;
        end else if(par_reset1_out) begin
            par_reset1_write_en = 1'd1;
        end else par_reset1_write_en = 1'd0;
        par_reset10_clk = clk;
        if(((par_done_reg25_out & par_done_reg26_out) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            par_reset10_in = 1'd1;
        end else if(par_reset10_out) begin
            par_reset10_in = 1'd0;
        end else par_reset10_in = 1'd0;
        if(((par_done_reg25_out & par_done_reg26_out) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            par_reset10_write_en = 1'd1;
        end else if(par_reset10_out) begin
            par_reset10_write_en = 1'd1;
        end else par_reset10_write_en = 1'd0;
        par_reset11_clk = clk;
        if(((par_done_reg27_out & par_done_reg28_out) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset11_in = 1'd1;
        end else if(par_reset11_out) begin
            par_reset11_in = 1'd0;
        end else par_reset11_in = 1'd0;
        if(((par_done_reg27_out & par_done_reg28_out) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset11_write_en = 1'd1;
        end else if(par_reset11_out) begin
            par_reset11_write_en = 1'd1;
        end else par_reset11_write_en = 1'd0;
        par_reset12_clk = clk;
        if(((par_done_reg29_out & par_done_reg30_out) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset12_in = 1'd1;
        end else if(par_reset12_out) begin
            par_reset12_in = 1'd0;
        end else par_reset12_in = 1'd0;
        if(((par_done_reg29_out & par_done_reg30_out) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset12_write_en = 1'd1;
        end else if(par_reset12_out) begin
            par_reset12_write_en = 1'd1;
        end else par_reset12_write_en = 1'd0;
        par_reset13_clk = clk;
        if(((par_done_reg31_out & par_done_reg32_out) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset13_in = 1'd1;
        end else if(par_reset13_out) begin
            par_reset13_in = 1'd0;
        end else par_reset13_in = 1'd0;
        if(((par_done_reg31_out & par_done_reg32_out) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset13_write_en = 1'd1;
        end else if(par_reset13_out) begin
            par_reset13_write_en = 1'd1;
        end else par_reset13_write_en = 1'd0;
        par_reset14_clk = clk;
        if(((par_done_reg33_out & par_done_reg34_out) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset14_in = 1'd1;
        end else if(par_reset14_out) begin
            par_reset14_in = 1'd0;
        end else par_reset14_in = 1'd0;
        if(((par_done_reg33_out & par_done_reg34_out) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset14_write_en = 1'd1;
        end else if(par_reset14_out) begin
            par_reset14_write_en = 1'd1;
        end else par_reset14_write_en = 1'd0;
        par_reset15_clk = clk;
        if(((par_done_reg35_out & par_done_reg36_out) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset15_in = 1'd1;
        end else if(par_reset15_out) begin
            par_reset15_in = 1'd0;
        end else par_reset15_in = 1'd0;
        if(((par_done_reg35_out & par_done_reg36_out) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset15_write_en = 1'd1;
        end else if(par_reset15_out) begin
            par_reset15_write_en = 1'd1;
        end else par_reset15_write_en = 1'd0;
        par_reset16_clk = clk;
        if(((par_done_reg37_out & par_done_reg38_out) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset16_in = 1'd1;
        end else if(par_reset16_out) begin
            par_reset16_in = 1'd0;
        end else par_reset16_in = 1'd0;
        if(((par_done_reg37_out & par_done_reg38_out) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset16_write_en = 1'd1;
        end else if(par_reset16_out) begin
            par_reset16_write_en = 1'd1;
        end else par_reset16_write_en = 1'd0;
        par_reset17_clk = clk;
        if(((par_done_reg39_out & par_done_reg40_out) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset17_in = 1'd1;
        end else if(par_reset17_out) begin
            par_reset17_in = 1'd0;
        end else par_reset17_in = 1'd0;
        if(((par_done_reg39_out & par_done_reg40_out) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset17_write_en = 1'd1;
        end else if(par_reset17_out) begin
            par_reset17_write_en = 1'd1;
        end else par_reset17_write_en = 1'd0;
        par_reset18_clk = clk;
        if(((par_done_reg41_out & par_done_reg42_out) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset18_in = 1'd1;
        end else if(par_reset18_out) begin
            par_reset18_in = 1'd0;
        end else par_reset18_in = 1'd0;
        if(((par_done_reg41_out & par_done_reg42_out) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            par_reset18_write_en = 1'd1;
        end else if(par_reset18_out) begin
            par_reset18_write_en = 1'd1;
        end else par_reset18_write_en = 1'd0;
        par_reset19_clk = clk;
        if(((par_done_reg43_out & par_done_reg44_out) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))) begin
            par_reset19_in = 1'd1;
        end else if(par_reset19_out) begin
            par_reset19_in = 1'd0;
        end else par_reset19_in = 1'd0;
        if(((par_done_reg43_out & par_done_reg44_out) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))) begin
            par_reset19_write_en = 1'd1;
        end else if(par_reset19_out) begin
            par_reset19_write_en = 1'd1;
        end else par_reset19_write_en = 1'd0;
        par_reset2_clk = clk;
        if(((par_done_reg5_out & par_done_reg6_out) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset2_in = 1'd1;
        end else if(par_reset2_out) begin
            par_reset2_in = 1'd0;
        end else par_reset2_in = 1'd0;
        if(((par_done_reg5_out & par_done_reg6_out) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset2_write_en = 1'd1;
        end else if(par_reset2_out) begin
            par_reset2_write_en = 1'd1;
        end else par_reset2_write_en = 1'd0;
        par_reset3_clk = clk;
        if(((par_done_reg7_out & par_done_reg8_out) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset3_in = 1'd1;
        end else if(par_reset3_out) begin
            par_reset3_in = 1'd0;
        end else par_reset3_in = 1'd0;
        if(((par_done_reg7_out & par_done_reg8_out) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset3_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_reset3_write_en = 1'd1;
        end else par_reset3_write_en = 1'd0;
        par_reset4_clk = clk;
        if(((par_done_reg9_out & par_done_reg10_out) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset4_in = 1'd1;
        end else if(par_reset4_out) begin
            par_reset4_in = 1'd0;
        end else par_reset4_in = 1'd0;
        if(((par_done_reg9_out & par_done_reg10_out) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset4_write_en = 1'd1;
        end else if(par_reset4_out) begin
            par_reset4_write_en = 1'd1;
        end else par_reset4_write_en = 1'd0;
        par_reset5_clk = clk;
        if(((par_done_reg11_out & par_done_reg12_out) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset5_in = 1'd1;
        end else if(par_reset5_out) begin
            par_reset5_in = 1'd0;
        end else par_reset5_in = 1'd0;
        if(((par_done_reg11_out & par_done_reg12_out) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            par_reset5_write_en = 1'd1;
        end else if(par_reset5_out) begin
            par_reset5_write_en = 1'd1;
        end else par_reset5_write_en = 1'd0;
        par_reset6_clk = clk;
        if(((((par_done_reg13_out & par_done_reg14_out) & par_done_reg15_out) & par_done_reg16_out) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_reset6_in = 1'd1;
        end else if(par_reset6_out) begin
            par_reset6_in = 1'd0;
        end else par_reset6_in = 1'd0;
        if(((((par_done_reg13_out & par_done_reg14_out) & par_done_reg15_out) & par_done_reg16_out) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))) begin
            par_reset6_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_reset6_write_en = 1'd1;
        end else par_reset6_write_en = 1'd0;
        par_reset7_clk = clk;
        if(((((par_done_reg17_out & par_done_reg18_out) & par_done_reg19_out) & par_done_reg20_out) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_reset7_in = 1'd1;
        end else if(par_reset7_out) begin
            par_reset7_in = 1'd0;
        end else par_reset7_in = 1'd0;
        if(((((par_done_reg17_out & par_done_reg18_out) & par_done_reg19_out) & par_done_reg20_out) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_reset7_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_reset7_write_en = 1'd1;
        end else par_reset7_write_en = 1'd0;
        par_reset8_clk = clk;
        if(((par_done_reg21_out & par_done_reg22_out) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_reset8_in = 1'd1;
        end else if(par_reset8_out) begin
            par_reset8_in = 1'd0;
        end else par_reset8_in = 1'd0;
        if(((par_done_reg21_out & par_done_reg22_out) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            par_reset8_write_en = 1'd1;
        end else if(par_reset8_out) begin
            par_reset8_write_en = 1'd1;
        end else par_reset8_write_en = 1'd0;
        par_reset9_clk = clk;
        if(((par_done_reg23_out & par_done_reg24_out) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            par_reset9_in = 1'd1;
        end else if(par_reset9_out) begin
            par_reset9_in = 1'd0;
        end else par_reset9_in = 1'd0;
        if(((par_done_reg23_out & par_done_reg24_out) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            par_reset9_write_en = 1'd1;
        end else if(par_reset9_out) begin
            par_reset9_write_en = 1'd1;
        end else par_reset9_write_en = 1'd0;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            rsh0_left = j0_out;
        end else if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            rsh0_left = j4_out;
        end else rsh0_left = 7'd0;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            rsh0_right = const10_out;
        end else if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            rsh0_right = const10_out;
        end else rsh0_right = 7'd0;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            rsh1_left = i1_out;
        end else if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            rsh1_left = i7_out;
        end else rsh1_left = 7'd0;
        if((((fsm1_out == 32'd1) & ~A0_0_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm1_out == 32'd3)) & (((fsm2_out == 32'd1) & ~done_reg0_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm2_out == 32'd3)) & (((fsm3_out == 32'd1) & ~done_reg1_out) & (~(par_done_reg16_out | (fsm3_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))))) begin
            rsh1_right = const11_out;
        end else if((((fsm14_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored10_out & cond_computed10_out) & ~(fsm14_out == 32'd3)) & (((fsm15_out == 32'd1) & ~done_reg10_out) & (((cond_stored11_out & cond_computed11_out) & ~(fsm15_out == 32'd3)) & (((fsm16_out == 32'd1) & ~done_reg11_out) & (~(par_done_reg44_out | (fsm16_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))))) begin
            rsh1_right = const11_out;
        end else rsh1_right = 7'd0;
        if((~(par_done_reg7_out | w0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else if((~(par_done_reg9_out | x0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else if((~(par_done_reg11_out | y0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else if((((fsm_out == 32'd8) & ~z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            rsh10_left = i0_out;
        end else if((~(par_done_reg_out | u10_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else if((((fsm12_out == 32'd0) & ~u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg30_out | v1_sh_read0_0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg32_out | u2_sh_read0_0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg1_out | v10_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else if((~(par_done_reg34_out | v2_sh_read0_0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg36_out | w_sh_read0_0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg38_out | x_sh_read0_0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg40_out | y_sh_read0_0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg42_out | z_sh_read0_0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_left = i6_out;
        end else if((~(par_done_reg3_out | u20_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else if((~(par_done_reg5_out | v20_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_left = i0_out;
        end else rsh10_left = 7'd0;
        if((~(par_done_reg7_out | w0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg9_out | x0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg11_out | y0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((((fsm_out == 32'd8) & ~z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg_out | u10_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((((fsm12_out == 32'd0) & ~u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg30_out | v1_sh_read0_0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg32_out | u2_sh_read0_0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg1_out | v10_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg34_out | v2_sh_read0_0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg36_out | w_sh_read0_0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg38_out | x_sh_read0_0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg40_out | y_sh_read0_0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg42_out | z_sh_read0_0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg3_out | u20_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else if((~(par_done_reg5_out | v20_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            rsh10_right = const13_out;
        end else rsh10_right = 7'd0;
        tmp1_0_clk = clk;
        if((((fsm4_out == 32'd2) & ~tmp1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            tmp1_0_in = add10_out;
        end else tmp1_0_in = 32'd0;
        if((((fsm4_out == 32'd2) & ~tmp1_0_done) & (~(par_done_reg21_out | (fsm4_out == 32'd3)) & (((fsm5_out == 32'd1) & ~par_reset8_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go))))))))) begin
            tmp1_0_write_en = 1'd1;
        end else tmp1_0_write_en = 1'd0;
        tmp2_0_clk = clk;
        if((((fsm7_out == 32'd3) & ~tmp2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            tmp2_0_in = bin_read3_0_out;
        end else tmp2_0_in = 32'd0;
        if((((fsm7_out == 32'd3) & ~tmp2_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            tmp2_0_write_en = 1'd1;
        end else tmp2_0_write_en = 1'd0;
        tmp3_0_clk = clk;
        if((~(par_done_reg25_out | tmp3_0_done) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            tmp3_0_in = z0_read_data;
        end else tmp3_0_in = 32'd0;
        if((~(par_done_reg25_out | tmp3_0_done) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            tmp3_0_write_en = 1'd1;
        end else tmp3_0_write_en = 1'd0;
        tmp4_0_clk = clk;
        if((((fsm10_out == 32'd3) & ~tmp4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            tmp4_0_in = bin_read5_0_out;
        end else tmp4_0_in = 32'd0;
        if((((fsm10_out == 32'd3) & ~tmp4_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            tmp4_0_write_en = 1'd1;
        end else tmp4_0_write_en = 1'd0;
        if((~(par_done_reg17_out | u1_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            u10_addr0 = i2_out;
        end else if((~(par_done_reg_out | u10_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u10_addr0 = rsh10_out;
        end else if((((fsm12_out == 32'd0) & ~u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            u10_addr0 = rsh10_out;
        end else u10_addr0 = 7'd0;
        u10_clk = clk;
        if((~(par_done_reg_out | u10_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u10_write_data = u1_int_read0_0_out;
        end else u10_write_data = 32'd0;
        if((~(par_done_reg_out | u10_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u10_write_en = 1'd1;
        end else u10_write_en = 1'd0;
        u1_int_read0_0_clk = clk;
        if((((fsm_out == 32'd0) & ~u1_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            u1_int_read0_0_in = u1_int0_read_data;
        end else u1_int_read0_0_in = 32'd0;
        if((((fsm_out == 32'd0) & ~u1_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            u1_int_read0_0_write_en = 1'd1;
        end else u1_int_read0_0_write_en = 1'd0;
        u1_read0_0_clk = clk;
        if((~(par_done_reg17_out | u1_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            u1_read0_0_in = u10_read_data;
        end else u1_read0_0_in = 32'd0;
        if((~(par_done_reg17_out | u1_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            u1_read0_0_write_en = 1'd1;
        end else u1_read0_0_write_en = 1'd0;
        u1_sh_read0_0_clk = clk;
        if((((fsm12_out == 32'd0) & ~u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            u1_sh_read0_0_in = u10_read_data;
        end else u1_sh_read0_0_in = 32'd0;
        if((((fsm12_out == 32'd0) & ~u1_sh_read0_0_done) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go))))))) begin
            u1_sh_read0_0_write_en = 1'd1;
        end else u1_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg19_out | u2_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            u20_addr0 = i2_out;
        end else if((~(par_done_reg32_out | u2_sh_read0_0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u20_addr0 = rsh10_out;
        end else if((~(par_done_reg3_out | u20_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u20_addr0 = rsh10_out;
        end else u20_addr0 = 7'd0;
        u20_clk = clk;
        if((~(par_done_reg3_out | u20_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u20_write_data = u2_int_read0_0_out;
        end else u20_write_data = 32'd0;
        if((~(par_done_reg3_out | u20_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u20_write_en = 1'd1;
        end else u20_write_en = 1'd0;
        u2_int_read0_0_clk = clk;
        if((~(par_done_reg2_out | u2_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u2_int_read0_0_in = u2_int0_read_data;
        end else u2_int_read0_0_in = 32'd0;
        if((~(par_done_reg2_out | u2_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            u2_int_read0_0_write_en = 1'd1;
        end else u2_int_read0_0_write_en = 1'd0;
        u2_read0_0_clk = clk;
        if((~(par_done_reg19_out | u2_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            u2_read0_0_in = u20_read_data;
        end else u2_read0_0_in = 32'd0;
        if((~(par_done_reg19_out | u2_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            u2_read0_0_write_en = 1'd1;
        end else u2_read0_0_write_en = 1'd0;
        u2_sh_read0_0_clk = clk;
        if((~(par_done_reg32_out | u2_sh_read0_0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u2_sh_read0_0_in = u20_read_data;
        end else u2_sh_read0_0_in = 32'd0;
        if((~(par_done_reg32_out | u2_sh_read0_0_done) & (((fsm12_out == 32'd2) & ~par_reset13_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            u2_sh_read0_0_write_en = 1'd1;
        end else u2_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg18_out | v1_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            v10_addr0 = j1_out;
        end else if((~(par_done_reg30_out | v1_sh_read0_0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v10_addr0 = rsh10_out;
        end else if((~(par_done_reg1_out | v10_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v10_addr0 = rsh10_out;
        end else v10_addr0 = 7'd0;
        v10_clk = clk;
        if((~(par_done_reg1_out | v10_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v10_write_data = v1_int_read0_0_out;
        end else v10_write_data = 32'd0;
        if((~(par_done_reg1_out | v10_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v10_write_en = 1'd1;
        end else v10_write_en = 1'd0;
        v1_int_read0_0_clk = clk;
        if((~(par_done_reg0_out | v1_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v1_int_read0_0_in = v1_int0_read_data;
        end else v1_int_read0_0_in = 32'd0;
        if((~(par_done_reg0_out | v1_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v1_int_read0_0_write_en = 1'd1;
        end else v1_int_read0_0_write_en = 1'd0;
        v1_read0_0_clk = clk;
        if((~(par_done_reg18_out | v1_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            v1_read0_0_in = v10_read_data;
        end else v1_read0_0_in = 32'd0;
        if((~(par_done_reg18_out | v1_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            v1_read0_0_write_en = 1'd1;
        end else v1_read0_0_write_en = 1'd0;
        v1_sh_read0_0_clk = clk;
        if((~(par_done_reg30_out | v1_sh_read0_0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v1_sh_read0_0_in = v10_read_data;
        end else v1_sh_read0_0_in = 32'd0;
        if((~(par_done_reg30_out | v1_sh_read0_0_done) & (((fsm12_out == 32'd1) & ~par_reset12_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v1_sh_read0_0_write_en = 1'd1;
        end else v1_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg20_out | v2_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            v20_addr0 = j1_out;
        end else if((~(par_done_reg34_out | v2_sh_read0_0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v20_addr0 = rsh10_out;
        end else if((~(par_done_reg5_out | v20_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v20_addr0 = rsh10_out;
        end else v20_addr0 = 7'd0;
        v20_clk = clk;
        if((~(par_done_reg5_out | v20_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v20_write_data = v2_int_read0_0_out;
        end else v20_write_data = 32'd0;
        if((~(par_done_reg5_out | v20_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v20_write_en = 1'd1;
        end else v20_write_en = 1'd0;
        v2_int_read0_0_clk = clk;
        if((~(par_done_reg4_out | v2_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v2_int_read0_0_in = v2_int0_read_data;
        end else v2_int_read0_0_in = 32'd0;
        if((~(par_done_reg4_out | v2_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            v2_int_read0_0_write_en = 1'd1;
        end else v2_int_read0_0_write_en = 1'd0;
        v2_read0_0_clk = clk;
        if((~(par_done_reg20_out | v2_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            v2_read0_0_in = v20_read_data;
        end else v2_read0_0_in = 32'd0;
        if((~(par_done_reg20_out | v2_read0_0_done) & (((fsm5_out == 32'd0) & ~par_reset7_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm5_out == 32'd4)) & (((fsm6_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm6_out == 32'd3)) & (((fsm17_out == 32'd2) & ~done_reg3_out) & (go | go)))))))) begin
            v2_read0_0_write_en = 1'd1;
        end else v2_read0_0_write_en = 1'd0;
        v2_sh_read0_0_clk = clk;
        if((~(par_done_reg34_out | v2_sh_read0_0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v2_sh_read0_0_in = v20_read_data;
        end else v2_sh_read0_0_in = 32'd0;
        if((~(par_done_reg34_out | v2_sh_read0_0_done) & (((fsm12_out == 32'd3) & ~par_reset14_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            v2_sh_read0_0_write_en = 1'd1;
        end else v2_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg7_out | w0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            w0_addr0 = rsh10_out;
        end else if((((fsm10_out == 32'd4) & ~w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            w0_addr0 = i5_out;
        end else if((((fsm10_out == 32'd4) & ~w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            w0_addr0 = i5_out;
        end else if((~(par_done_reg36_out | w_sh_read0_0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            w0_addr0 = rsh10_out;
        end else w0_addr0 = 7'd0;
        w0_clk = clk;
        if((~(par_done_reg7_out | w0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            w0_write_data = w_int_read0_0_out;
        end else if((((fsm10_out == 32'd4) & ~w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            w0_write_data = add10_out;
        end else w0_write_data = 32'd0;
        if((~(par_done_reg7_out | w0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            w0_write_en = 1'd1;
        end else if((((fsm10_out == 32'd4) & ~w0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go))))))) begin
            w0_write_en = 1'd1;
        end else w0_write_en = 1'd0;
        w_int_read0_0_clk = clk;
        if((~(par_done_reg6_out | w_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            w_int_read0_0_in = w_int0_read_data;
        end else w_int_read0_0_in = 32'd0;
        if((~(par_done_reg6_out | w_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            w_int_read0_0_write_en = 1'd1;
        end else w_int_read0_0_write_en = 1'd0;
        w_sh_read0_0_clk = clk;
        if((~(par_done_reg36_out | w_sh_read0_0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            w_sh_read0_0_in = w0_read_data;
        end else w_sh_read0_0_in = 32'd0;
        if((~(par_done_reg36_out | w_sh_read0_0_done) & (((fsm12_out == 32'd4) & ~par_reset15_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            w_sh_read0_0_write_en = 1'd1;
        end else w_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg9_out | x0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            x0_addr0 = rsh10_out;
        end else if((((fsm7_out == 32'd4) & ~x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            x0_addr0 = i3_out;
        end else if((((fsm7_out == 32'd4) & ~x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            x0_addr0 = i3_out;
        end else if((~(par_done_reg26_out | old_1_done) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            x0_addr0 = i4_out;
        end else if((((fsm9_out == 32'd1) & ~x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            x0_addr0 = i4_out;
        end else if((~(par_done_reg28_out | x_read0_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            x0_addr0 = j3_out;
        end else if((~(par_done_reg38_out | x_sh_read0_0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            x0_addr0 = rsh10_out;
        end else x0_addr0 = 7'd0;
        x0_clk = clk;
        if((~(par_done_reg9_out | x0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            x0_write_data = x_int_read0_0_out;
        end else if((((fsm7_out == 32'd4) & ~x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            x0_write_data = add10_out;
        end else if((((fsm9_out == 32'd1) & ~x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            x0_write_data = add10_out;
        end else x0_write_data = 32'd0;
        if((~(par_done_reg9_out | x0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            x0_write_en = 1'd1;
        end else if((((fsm7_out == 32'd4) & ~x0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go))))))) begin
            x0_write_en = 1'd1;
        end else if((((fsm9_out == 32'd1) & ~x0_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go))))) begin
            x0_write_en = 1'd1;
        end else x0_write_en = 1'd0;
        x_int_read0_0_clk = clk;
        if((~(par_done_reg8_out | x_int_read0_0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            x_int_read0_0_in = x_int0_read_data;
        end else x_int_read0_0_in = 32'd0;
        if((~(par_done_reg8_out | x_int_read0_0_done) & (((fsm_out == 32'd5) & ~par_reset3_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            x_int_read0_0_write_en = 1'd1;
        end else x_int_read0_0_write_en = 1'd0;
        x_read0_0_clk = clk;
        if((~(par_done_reg28_out | x_read0_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            x_read0_0_in = x0_read_data;
        end else x_read0_0_in = 32'd0;
        if((~(par_done_reg28_out | x_read0_0_done) & (((fsm10_out == 32'd0) & ~par_reset11_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm10_out == 32'd6)) & (((fsm11_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm11_out == 32'd3)) & (((fsm17_out == 32'd8) & ~done_reg8_out) & (go | go)))))))) begin
            x_read0_0_write_en = 1'd1;
        end else x_read0_0_write_en = 1'd0;
        x_sh_read0_0_clk = clk;
        if((~(par_done_reg38_out | x_sh_read0_0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            x_sh_read0_0_in = x0_read_data;
        end else x_sh_read0_0_in = 32'd0;
        if((~(par_done_reg38_out | x_sh_read0_0_done) & (((fsm12_out == 32'd5) & ~par_reset16_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            x_sh_read0_0_write_en = 1'd1;
        end else x_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg11_out | y0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            y0_addr0 = rsh10_out;
        end else if((~(par_done_reg24_out | y_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            y0_addr0 = j2_out;
        end else if((~(par_done_reg40_out | y_sh_read0_0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            y0_addr0 = rsh10_out;
        end else y0_addr0 = 7'd0;
        y0_clk = clk;
        if((~(par_done_reg11_out | y0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            y0_write_data = y_int_read0_0_out;
        end else y0_write_data = 32'd0;
        if((~(par_done_reg11_out | y0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            y0_write_en = 1'd1;
        end else y0_write_en = 1'd0;
        y_int_read0_0_clk = clk;
        if((~(par_done_reg10_out | y_int_read0_0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            y_int_read0_0_in = y_int0_read_data;
        end else y_int_read0_0_in = 32'd0;
        if((~(par_done_reg10_out | y_int_read0_0_done) & (((fsm_out == 32'd6) & ~par_reset4_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            y_int_read0_0_write_en = 1'd1;
        end else y_int_read0_0_write_en = 1'd0;
        y_read0_0_clk = clk;
        if((~(par_done_reg24_out | y_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            y_read0_0_in = y0_read_data;
        end else y_read0_0_in = 32'd0;
        if((~(par_done_reg24_out | y_read0_0_done) & (((fsm7_out == 32'd0) & ~par_reset9_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm7_out == 32'd6)) & (((fsm8_out == 32'd1) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm8_out == 32'd3)) & (((fsm17_out == 32'd4) & ~done_reg5_out) & (go | go)))))))) begin
            y_read0_0_write_en = 1'd1;
        end else y_read0_0_write_en = 1'd0;
        y_sh_read0_0_clk = clk;
        if((~(par_done_reg40_out | y_sh_read0_0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            y_sh_read0_0_in = y0_read_data;
        end else y_sh_read0_0_in = 32'd0;
        if((~(par_done_reg40_out | y_sh_read0_0_done) & (((fsm12_out == 32'd6) & ~par_reset17_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            y_sh_read0_0_write_en = 1'd1;
        end else y_sh_read0_0_write_en = 1'd0;
        if((((fsm_out == 32'd8) & ~z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            z0_addr0 = rsh10_out;
        end else if((~(par_done_reg25_out | tmp3_0_done) & (((fsm9_out == 32'd0) & ~par_reset10_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm9_out == 32'd3)) & (((fsm17_out == 32'd6) & ~done_reg6_out) & (go | go)))))) begin
            z0_addr0 = i4_out;
        end else if((~(par_done_reg42_out | z_sh_read0_0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            z0_addr0 = rsh10_out;
        end else z0_addr0 = 7'd0;
        z0_clk = clk;
        if((((fsm_out == 32'd8) & ~z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            z0_write_data = z_int_read0_0_out;
        end else z0_write_data = 32'd0;
        if((((fsm_out == 32'd8) & ~z0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go))))))) begin
            z0_write_en = 1'd1;
        end else z0_write_en = 1'd0;
        z_int_read0_0_clk = clk;
        if((~(par_done_reg12_out | z_int_read0_0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            z_int_read0_0_in = z_int0_read_data;
        end else z_int_read0_0_in = 32'd0;
        if((~(par_done_reg12_out | z_int_read0_0_done) & (((fsm_out == 32'd7) & ~par_reset5_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd10)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (~(par_done_reg15_out | (fsm0_out == 32'd2)) & (((fsm17_out == 32'd0) & ~par_reset6_out) & (go | go)))))))) begin
            z_int_read0_0_write_en = 1'd1;
        end else z_int_read0_0_write_en = 1'd0;
        z_sh_read0_0_clk = clk;
        if((~(par_done_reg42_out | z_sh_read0_0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            z_sh_read0_0_in = z0_read_data;
        end else z_sh_read0_0_in = 32'd0;
        if((~(par_done_reg42_out | z_sh_read0_0_done) & (((fsm12_out == 32'd7) & ~par_reset18_out) & (((cond_stored9_out & cond_computed9_out) & ~(fsm12_out == 32'd10)) & (((fsm13_out == 32'd1) & ~done_reg9_out) & (~(par_done_reg43_out | (fsm13_out == 32'd2)) & (((fsm17_out == 32'd9) & ~par_reset19_out) & (go | go)))))))) begin
            z_sh_read0_0_write_en = 1'd1;
        end else z_sh_read0_0_write_en = 1'd0;
    end
endmodule
