module std_add
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left + right;
endmodule
module std_const
  #(parameter width = 32,
    parameter value = 0)
   (output logic [width - 1:0] out);
  assign out = value;
endmodule
module std_le
  #(parameter width = 32)
  (input logic [width-1:0] left,
   input logic [width-1:0] right,
   output logic            out);
  assign out = left <= right;
endmodule
module std_mem_d2
  #(parameter width = 32,
    parameter d0_size = 16,
    parameter d1_size = 16,
    parameter d0_idx_size = 4,
    parameter d1_idx_size = 4)
   (input logic [d0_idx_size-1:0] addr0,
    input logic [d1_idx_size-1:0] addr1,
    input logic [width-1:0]   write_data,
    input logic               write_en,
    input logic               clk,
    output logic [width-1:0]  read_data,
    output logic done);

  /* verilator lint_off WIDTH */
  logic [width-1:0]  mem[d0_size-1:0][d1_size-1:0];

  assign read_data = mem[addr0][addr1];
  always_ff @(posedge clk) begin
    if (write_en) begin
      mem[addr0][addr1] <= write_data;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule
module std_mult_pipe
  #(parameter width = 32)
   (input logic [width-1:0] left,
    input logic [width-1:0] right,
    input logic go,
    input logic clk,
    output logic [width-1:0] out,
    output logic done);
   logic [width-1:0] rtmp;
   logic [width-1:0] ltmp;
   logic [width-1:0] out_tmp;
   reg done_buf[1:0];
   always_ff @(posedge clk) begin
     if (go) begin
       rtmp <= right;
       ltmp <= left;
       out_tmp <= rtmp * ltmp;
       out <= out_tmp;

       done <= done_buf[1];
       done_buf[0] <= 1'b1;
       done_buf[1] <= done_buf[0];
     end else begin
       rtmp <= 0;
       ltmp <= 0;
       out_tmp <= 0;
       out <= 0;

       done <= 0;
       done_buf[0] <= 0;
       done_buf[1] <= 0;
     end
   end
 endmodule
module std_reg
  #(parameter width = 32)
   (input wire [width-1:0] in,
    input wire write_en,
    input wire clk,
    // output
    output logic [width - 1:0] out,
    output logic done);

  always_ff @(posedge clk) begin
    if (write_en) begin
      out <= in;
      done <= 1'd1;
    end else
      done <= 1'd0;
  end
endmodule
module std_rsh
  #(parameter width = 32)
  (input  logic [width-1:0] left,
    input  logic [width-1:0] right,
    output logic [width-1:0] out);
  assign out = left >> right;
endmodule
module main (
    input logic go,
    input logic clk,
    output logic done,
    output logic [3:0] A_int0_0_addr0,
    output logic [3:0] A_int0_0_addr1,
    output logic [31:0] A_int0_0_write_data,
    output logic A_int0_0_write_en,
    output logic A_int0_0_clk,
    input logic [31:0] A_int0_0_read_data,
    input logic A_int0_0_done,
    output logic [3:0] B_int0_0_addr0,
    output logic [3:0] B_int0_0_addr1,
    output logic [31:0] B_int0_0_write_data,
    output logic B_int0_0_write_en,
    output logic B_int0_0_clk,
    input logic [31:0] B_int0_0_read_data,
    input logic B_int0_0_done,
    output logic [3:0] C_int0_0_addr0,
    output logic [3:0] C_int0_0_addr1,
    output logic [31:0] C_int0_0_write_data,
    output logic C_int0_0_write_en,
    output logic C_int0_0_clk,
    input logic [31:0] C_int0_0_read_data,
    input logic C_int0_0_done,
    output logic [3:0] D_int0_0_addr0,
    output logic [3:0] D_int0_0_addr1,
    output logic [31:0] D_int0_0_write_data,
    output logic D_int0_0_write_en,
    output logic D_int0_0_clk,
    input logic [31:0] D_int0_0_read_data,
    input logic D_int0_0_done,
    output logic alpha_int0_addr0,
    output logic [31:0] alpha_int0_write_data,
    output logic alpha_int0_write_en,
    output logic alpha_int0_clk,
    input logic [31:0] alpha_int0_read_data,
    input logic alpha_int0_done,
    output logic beta_int0_addr0,
    output logic [31:0] beta_int0_write_data,
    output logic beta_int0_write_en,
    output logic beta_int0_clk,
    input logic [31:0] beta_int0_read_data,
    input logic beta_int0_done,
    output logic [3:0] tmp_int0_0_addr0,
    output logic [3:0] tmp_int0_0_addr1,
    output logic [31:0] tmp_int0_0_write_data,
    output logic tmp_int0_0_write_en,
    output logic tmp_int0_0_clk,
    input logic [31:0] tmp_int0_0_read_data,
    input logic tmp_int0_0_done
);
    logic [3:0] A0_0_addr0;
    logic [3:0] A0_0_addr1;
    logic [31:0] A0_0_write_data;
    logic A0_0_write_en;
    logic A0_0_clk;
    logic [31:0] A0_0_read_data;
    logic A0_0_done;
    logic [31:0] A_int_read0_0_in;
    logic A_int_read0_0_write_en;
    logic A_int_read0_0_clk;
    logic [31:0] A_int_read0_0_out;
    logic A_int_read0_0_done;
    logic [31:0] A_read0_0_in;
    logic A_read0_0_write_en;
    logic A_read0_0_clk;
    logic [31:0] A_read0_0_out;
    logic A_read0_0_done;
    logic [31:0] A_sh_read0_0_in;
    logic A_sh_read0_0_write_en;
    logic A_sh_read0_0_clk;
    logic [31:0] A_sh_read0_0_out;
    logic A_sh_read0_0_done;
    logic [3:0] B0_0_addr0;
    logic [3:0] B0_0_addr1;
    logic [31:0] B0_0_write_data;
    logic B0_0_write_en;
    logic B0_0_clk;
    logic [31:0] B0_0_read_data;
    logic B0_0_done;
    logic [31:0] B_int_read0_0_in;
    logic B_int_read0_0_write_en;
    logic B_int_read0_0_clk;
    logic [31:0] B_int_read0_0_out;
    logic B_int_read0_0_done;
    logic [31:0] B_read0_0_in;
    logic B_read0_0_write_en;
    logic B_read0_0_clk;
    logic [31:0] B_read0_0_out;
    logic B_read0_0_done;
    logic [31:0] B_sh_read0_0_in;
    logic B_sh_read0_0_write_en;
    logic B_sh_read0_0_clk;
    logic [31:0] B_sh_read0_0_out;
    logic B_sh_read0_0_done;
    logic [3:0] C0_0_addr0;
    logic [3:0] C0_0_addr1;
    logic [31:0] C0_0_write_data;
    logic C0_0_write_en;
    logic C0_0_clk;
    logic [31:0] C0_0_read_data;
    logic C0_0_done;
    logic [31:0] C_int_read0_0_in;
    logic C_int_read0_0_write_en;
    logic C_int_read0_0_clk;
    logic [31:0] C_int_read0_0_out;
    logic C_int_read0_0_done;
    logic [31:0] C_read0_0_in;
    logic C_read0_0_write_en;
    logic C_read0_0_clk;
    logic [31:0] C_read0_0_out;
    logic C_read0_0_done;
    logic [31:0] C_sh_read0_0_in;
    logic C_sh_read0_0_write_en;
    logic C_sh_read0_0_clk;
    logic [31:0] C_sh_read0_0_out;
    logic C_sh_read0_0_done;
    logic [3:0] D0_0_addr0;
    logic [3:0] D0_0_addr1;
    logic [31:0] D0_0_write_data;
    logic D0_0_write_en;
    logic D0_0_clk;
    logic [31:0] D0_0_read_data;
    logic D0_0_done;
    logic [31:0] D_int_read0_0_in;
    logic D_int_read0_0_write_en;
    logic D_int_read0_0_clk;
    logic [31:0] D_int_read0_0_out;
    logic D_int_read0_0_done;
    logic [31:0] D_sh_read0_0_in;
    logic D_sh_read0_0_write_en;
    logic D_sh_read0_0_clk;
    logic [31:0] D_sh_read0_0_out;
    logic D_sh_read0_0_done;
    logic [3:0] add0_left;
    logic [3:0] add0_right;
    logic [3:0] add0_out;
    logic [31:0] add2_left;
    logic [31:0] add2_right;
    logic [31:0] add2_out;
    logic [31:0] alpha_int_read0_0_in;
    logic alpha_int_read0_0_write_en;
    logic alpha_int_read0_0_clk;
    logic [31:0] alpha_int_read0_0_out;
    logic alpha_int_read0_0_done;
    logic [31:0] beta_int_read0_0_in;
    logic beta_int_read0_0_write_en;
    logic beta_int_read0_0_clk;
    logic [31:0] beta_int_read0_0_out;
    logic beta_int_read0_0_done;
    logic [31:0] bin_read0_0_in;
    logic bin_read0_0_write_en;
    logic bin_read0_0_clk;
    logic [31:0] bin_read0_0_out;
    logic bin_read0_0_done;
    logic [31:0] bin_read1_0_in;
    logic bin_read1_0_write_en;
    logic bin_read1_0_clk;
    logic [31:0] bin_read1_0_out;
    logic bin_read1_0_done;
    logic [31:0] bin_read2_0_in;
    logic bin_read2_0_write_en;
    logic bin_read2_0_clk;
    logic [31:0] bin_read2_0_out;
    logic bin_read2_0_done;
    logic [31:0] bin_read3_0_in;
    logic bin_read3_0_write_en;
    logic bin_read3_0_clk;
    logic [31:0] bin_read3_0_out;
    logic bin_read3_0_done;
    logic [3:0] const0_out;
    logic [3:0] const1_out;
    logic [3:0] const10_out;
    logic [3:0] const14_out;
    logic [31:0] const20_out;
    logic const23_out;
    logic [31:0] d_tmp_0_in;
    logic d_tmp_0_write_en;
    logic d_tmp_0_clk;
    logic [31:0] d_tmp_0_out;
    logic d_tmp_0_done;
    logic [3:0] i0_in;
    logic i0_write_en;
    logic i0_clk;
    logic [3:0] i0_out;
    logic i0_done;
    logic [3:0] i00_in;
    logic i00_write_en;
    logic i00_clk;
    logic [3:0] i00_out;
    logic i00_done;
    logic [3:0] i01_in;
    logic i01_write_en;
    logic i01_clk;
    logic [3:0] i01_out;
    logic i01_done;
    logic [3:0] i10_in;
    logic i10_write_en;
    logic i10_clk;
    logic [3:0] i10_out;
    logic i10_done;
    logic [3:0] j0_in;
    logic j0_write_en;
    logic j0_clk;
    logic [3:0] j0_out;
    logic j0_done;
    logic [3:0] j00_in;
    logic j00_write_en;
    logic j00_clk;
    logic [3:0] j00_out;
    logic j00_done;
    logic [3:0] j01_in;
    logic j01_write_en;
    logic j01_clk;
    logic [3:0] j01_out;
    logic j01_done;
    logic [3:0] j10_in;
    logic j10_write_en;
    logic j10_clk;
    logic [3:0] j10_out;
    logic j10_done;
    logic [3:0] k0_in;
    logic k0_write_en;
    logic k0_clk;
    logic [3:0] k0_out;
    logic k0_done;
    logic [3:0] k10_in;
    logic k10_write_en;
    logic k10_clk;
    logic [3:0] k10_out;
    logic k10_done;
    logic [3:0] le0_left;
    logic [3:0] le0_right;
    logic le0_out;
    logic [31:0] mult_pipe0_left;
    logic [31:0] mult_pipe0_right;
    logic mult_pipe0_go;
    logic mult_pipe0_clk;
    logic [31:0] mult_pipe0_out;
    logic mult_pipe0_done;
    logic [31:0] mult_pipe1_left;
    logic [31:0] mult_pipe1_right;
    logic mult_pipe1_go;
    logic mult_pipe1_clk;
    logic [31:0] mult_pipe1_out;
    logic mult_pipe1_done;
    logic [31:0] mult_pipe2_left;
    logic [31:0] mult_pipe2_right;
    logic mult_pipe2_go;
    logic mult_pipe2_clk;
    logic [31:0] mult_pipe2_out;
    logic mult_pipe2_done;
    logic [31:0] mult_pipe3_left;
    logic [31:0] mult_pipe3_right;
    logic mult_pipe3_go;
    logic mult_pipe3_clk;
    logic [31:0] mult_pipe3_out;
    logic mult_pipe3_done;
    logic [3:0] rsh0_left;
    logic [3:0] rsh0_right;
    logic [3:0] rsh0_out;
    logic [3:0] rsh1_left;
    logic [3:0] rsh1_right;
    logic [3:0] rsh1_out;
    logic [3:0] tmp0_0_addr0;
    logic [3:0] tmp0_0_addr1;
    logic [31:0] tmp0_0_write_data;
    logic tmp0_0_write_en;
    logic tmp0_0_clk;
    logic [31:0] tmp0_0_read_data;
    logic tmp0_0_done;
    logic [31:0] tmp_int_read0_0_in;
    logic tmp_int_read0_0_write_en;
    logic tmp_int_read0_0_clk;
    logic [31:0] tmp_int_read0_0_out;
    logic tmp_int_read0_0_done;
    logic [31:0] tmp_read0_0_in;
    logic tmp_read0_0_write_en;
    logic tmp_read0_0_clk;
    logic [31:0] tmp_read0_0_out;
    logic tmp_read0_0_done;
    logic [31:0] tmp_sh_read0_0_in;
    logic tmp_sh_read0_0_write_en;
    logic tmp_sh_read0_0_clk;
    logic [31:0] tmp_sh_read0_0_out;
    logic tmp_sh_read0_0_done;
    logic [31:0] v1_0_in;
    logic v1_0_write_en;
    logic v1_0_clk;
    logic [31:0] v1_0_out;
    logic v1_0_done;
    logic [31:0] v_0_in;
    logic v_0_write_en;
    logic v_0_clk;
    logic [31:0] v_0_out;
    logic v_0_done;
    logic par_reset_in;
    logic par_reset_write_en;
    logic par_reset_clk;
    logic par_reset_out;
    logic par_reset_done;
    logic par_done_reg_in;
    logic par_done_reg_write_en;
    logic par_done_reg_clk;
    logic par_done_reg_out;
    logic par_done_reg_done;
    logic par_done_reg0_in;
    logic par_done_reg0_write_en;
    logic par_done_reg0_clk;
    logic par_done_reg0_out;
    logic par_done_reg0_done;
    logic par_reset0_in;
    logic par_reset0_write_en;
    logic par_reset0_clk;
    logic par_reset0_out;
    logic par_reset0_done;
    logic par_done_reg1_in;
    logic par_done_reg1_write_en;
    logic par_done_reg1_clk;
    logic par_done_reg1_out;
    logic par_done_reg1_done;
    logic par_done_reg2_in;
    logic par_done_reg2_write_en;
    logic par_done_reg2_clk;
    logic par_done_reg2_out;
    logic par_done_reg2_done;
    logic par_reset1_in;
    logic par_reset1_write_en;
    logic par_reset1_clk;
    logic par_reset1_out;
    logic par_reset1_done;
    logic par_done_reg3_in;
    logic par_done_reg3_write_en;
    logic par_done_reg3_clk;
    logic par_done_reg3_out;
    logic par_done_reg3_done;
    logic par_done_reg4_in;
    logic par_done_reg4_write_en;
    logic par_done_reg4_clk;
    logic par_done_reg4_out;
    logic par_done_reg4_done;
    logic par_reset2_in;
    logic par_reset2_write_en;
    logic par_reset2_clk;
    logic par_reset2_out;
    logic par_reset2_done;
    logic par_done_reg5_in;
    logic par_done_reg5_write_en;
    logic par_done_reg5_clk;
    logic par_done_reg5_out;
    logic par_done_reg5_done;
    logic par_done_reg6_in;
    logic par_done_reg6_write_en;
    logic par_done_reg6_clk;
    logic par_done_reg6_out;
    logic par_done_reg6_done;
    logic [31:0] fsm_in;
    logic fsm_write_en;
    logic fsm_clk;
    logic [31:0] fsm_out;
    logic fsm_done;
    logic cond_computed_in;
    logic cond_computed_write_en;
    logic cond_computed_clk;
    logic cond_computed_out;
    logic cond_computed_done;
    logic cond_stored_in;
    logic cond_stored_write_en;
    logic cond_stored_clk;
    logic cond_stored_out;
    logic cond_stored_done;
    logic done_reg_in;
    logic done_reg_write_en;
    logic done_reg_clk;
    logic done_reg_out;
    logic done_reg_done;
    logic [31:0] fsm0_in;
    logic fsm0_write_en;
    logic fsm0_clk;
    logic [31:0] fsm0_out;
    logic fsm0_done;
    logic cond_computed0_in;
    logic cond_computed0_write_en;
    logic cond_computed0_clk;
    logic cond_computed0_out;
    logic cond_computed0_done;
    logic cond_stored0_in;
    logic cond_stored0_write_en;
    logic cond_stored0_clk;
    logic cond_stored0_out;
    logic cond_stored0_done;
    logic done_reg0_in;
    logic done_reg0_write_en;
    logic done_reg0_clk;
    logic done_reg0_out;
    logic done_reg0_done;
    logic par_reset3_in;
    logic par_reset3_write_en;
    logic par_reset3_clk;
    logic par_reset3_out;
    logic par_reset3_done;
    logic par_done_reg7_in;
    logic par_done_reg7_write_en;
    logic par_done_reg7_clk;
    logic par_done_reg7_out;
    logic par_done_reg7_done;
    logic par_done_reg8_in;
    logic par_done_reg8_write_en;
    logic par_done_reg8_clk;
    logic par_done_reg8_out;
    logic par_done_reg8_done;
    logic par_done_reg9_in;
    logic par_done_reg9_write_en;
    logic par_done_reg9_clk;
    logic par_done_reg9_out;
    logic par_done_reg9_done;
    logic [31:0] fsm1_in;
    logic fsm1_write_en;
    logic fsm1_clk;
    logic [31:0] fsm1_out;
    logic fsm1_done;
    logic cond_computed1_in;
    logic cond_computed1_write_en;
    logic cond_computed1_clk;
    logic cond_computed1_out;
    logic cond_computed1_done;
    logic cond_stored1_in;
    logic cond_stored1_write_en;
    logic cond_stored1_clk;
    logic cond_stored1_out;
    logic cond_stored1_done;
    logic done_reg1_in;
    logic done_reg1_write_en;
    logic done_reg1_clk;
    logic done_reg1_out;
    logic done_reg1_done;
    logic [31:0] fsm2_in;
    logic fsm2_write_en;
    logic fsm2_clk;
    logic [31:0] fsm2_out;
    logic fsm2_done;
    logic cond_computed2_in;
    logic cond_computed2_write_en;
    logic cond_computed2_clk;
    logic cond_computed2_out;
    logic cond_computed2_done;
    logic cond_stored2_in;
    logic cond_stored2_write_en;
    logic cond_stored2_clk;
    logic cond_stored2_out;
    logic cond_stored2_done;
    logic done_reg2_in;
    logic done_reg2_write_en;
    logic done_reg2_clk;
    logic done_reg2_out;
    logic done_reg2_done;
    logic [31:0] fsm3_in;
    logic fsm3_write_en;
    logic fsm3_clk;
    logic [31:0] fsm3_out;
    logic fsm3_done;
    logic cond_computed3_in;
    logic cond_computed3_write_en;
    logic cond_computed3_clk;
    logic cond_computed3_out;
    logic cond_computed3_done;
    logic cond_stored3_in;
    logic cond_stored3_write_en;
    logic cond_stored3_clk;
    logic cond_stored3_out;
    logic cond_stored3_done;
    logic done_reg3_in;
    logic done_reg3_write_en;
    logic done_reg3_clk;
    logic done_reg3_out;
    logic done_reg3_done;
    logic par_reset4_in;
    logic par_reset4_write_en;
    logic par_reset4_clk;
    logic par_reset4_out;
    logic par_reset4_done;
    logic par_done_reg10_in;
    logic par_done_reg10_write_en;
    logic par_done_reg10_clk;
    logic par_done_reg10_out;
    logic par_done_reg10_done;
    logic par_done_reg11_in;
    logic par_done_reg11_write_en;
    logic par_done_reg11_clk;
    logic par_done_reg11_out;
    logic par_done_reg11_done;
    logic [31:0] fsm4_in;
    logic fsm4_write_en;
    logic fsm4_clk;
    logic [31:0] fsm4_out;
    logic fsm4_done;
    logic cond_computed4_in;
    logic cond_computed4_write_en;
    logic cond_computed4_clk;
    logic cond_computed4_out;
    logic cond_computed4_done;
    logic cond_stored4_in;
    logic cond_stored4_write_en;
    logic cond_stored4_clk;
    logic cond_stored4_out;
    logic cond_stored4_done;
    logic done_reg4_in;
    logic done_reg4_write_en;
    logic done_reg4_clk;
    logic done_reg4_out;
    logic done_reg4_done;
    logic [31:0] fsm5_in;
    logic fsm5_write_en;
    logic fsm5_clk;
    logic [31:0] fsm5_out;
    logic fsm5_done;
    logic cond_computed5_in;
    logic cond_computed5_write_en;
    logic cond_computed5_clk;
    logic cond_computed5_out;
    logic cond_computed5_done;
    logic cond_stored5_in;
    logic cond_stored5_write_en;
    logic cond_stored5_clk;
    logic cond_stored5_out;
    logic cond_stored5_done;
    logic done_reg5_in;
    logic done_reg5_write_en;
    logic done_reg5_clk;
    logic done_reg5_out;
    logic done_reg5_done;
    logic [31:0] fsm6_in;
    logic fsm6_write_en;
    logic fsm6_clk;
    logic [31:0] fsm6_out;
    logic fsm6_done;
    logic cond_computed6_in;
    logic cond_computed6_write_en;
    logic cond_computed6_clk;
    logic cond_computed6_out;
    logic cond_computed6_done;
    logic cond_stored6_in;
    logic cond_stored6_write_en;
    logic cond_stored6_clk;
    logic cond_stored6_out;
    logic cond_stored6_done;
    logic done_reg6_in;
    logic done_reg6_write_en;
    logic done_reg6_clk;
    logic done_reg6_out;
    logic done_reg6_done;
    logic par_reset5_in;
    logic par_reset5_write_en;
    logic par_reset5_clk;
    logic par_reset5_out;
    logic par_reset5_done;
    logic par_done_reg12_in;
    logic par_done_reg12_write_en;
    logic par_done_reg12_clk;
    logic par_done_reg12_out;
    logic par_done_reg12_done;
    logic par_done_reg13_in;
    logic par_done_reg13_write_en;
    logic par_done_reg13_clk;
    logic par_done_reg13_out;
    logic par_done_reg13_done;
    logic par_reset6_in;
    logic par_reset6_write_en;
    logic par_reset6_clk;
    logic par_reset6_out;
    logic par_reset6_done;
    logic par_done_reg14_in;
    logic par_done_reg14_write_en;
    logic par_done_reg14_clk;
    logic par_done_reg14_out;
    logic par_done_reg14_done;
    logic par_done_reg15_in;
    logic par_done_reg15_write_en;
    logic par_done_reg15_clk;
    logic par_done_reg15_out;
    logic par_done_reg15_done;
    logic par_reset7_in;
    logic par_reset7_write_en;
    logic par_reset7_clk;
    logic par_reset7_out;
    logic par_reset7_done;
    logic par_done_reg16_in;
    logic par_done_reg16_write_en;
    logic par_done_reg16_clk;
    logic par_done_reg16_out;
    logic par_done_reg16_done;
    logic par_done_reg17_in;
    logic par_done_reg17_write_en;
    logic par_done_reg17_clk;
    logic par_done_reg17_out;
    logic par_done_reg17_done;
    logic par_reset8_in;
    logic par_reset8_write_en;
    logic par_reset8_clk;
    logic par_reset8_out;
    logic par_reset8_done;
    logic par_done_reg18_in;
    logic par_done_reg18_write_en;
    logic par_done_reg18_clk;
    logic par_done_reg18_out;
    logic par_done_reg18_done;
    logic par_done_reg19_in;
    logic par_done_reg19_write_en;
    logic par_done_reg19_clk;
    logic par_done_reg19_out;
    logic par_done_reg19_done;
    logic [31:0] fsm7_in;
    logic fsm7_write_en;
    logic fsm7_clk;
    logic [31:0] fsm7_out;
    logic fsm7_done;
    logic cond_computed7_in;
    logic cond_computed7_write_en;
    logic cond_computed7_clk;
    logic cond_computed7_out;
    logic cond_computed7_done;
    logic cond_stored7_in;
    logic cond_stored7_write_en;
    logic cond_stored7_clk;
    logic cond_stored7_out;
    logic cond_stored7_done;
    logic done_reg7_in;
    logic done_reg7_write_en;
    logic done_reg7_clk;
    logic done_reg7_out;
    logic done_reg7_done;
    logic [31:0] fsm8_in;
    logic fsm8_write_en;
    logic fsm8_clk;
    logic [31:0] fsm8_out;
    logic fsm8_done;
    logic cond_computed8_in;
    logic cond_computed8_write_en;
    logic cond_computed8_clk;
    logic cond_computed8_out;
    logic cond_computed8_done;
    logic cond_stored8_in;
    logic cond_stored8_write_en;
    logic cond_stored8_clk;
    logic cond_stored8_out;
    logic cond_stored8_done;
    logic done_reg8_in;
    logic done_reg8_write_en;
    logic done_reg8_clk;
    logic done_reg8_out;
    logic done_reg8_done;
    logic [31:0] fsm9_in;
    logic fsm9_write_en;
    logic fsm9_clk;
    logic [31:0] fsm9_out;
    logic fsm9_done;
    initial begin
        A0_0_addr0 = 4'd0;
        A0_0_addr1 = 4'd0;
        A0_0_write_data = 32'd0;
        A0_0_write_en = 1'd0;
        A0_0_clk = 1'd0;
        A_int_read0_0_in = 32'd0;
        A_int_read0_0_write_en = 1'd0;
        A_int_read0_0_clk = 1'd0;
        A_read0_0_in = 32'd0;
        A_read0_0_write_en = 1'd0;
        A_read0_0_clk = 1'd0;
        A_sh_read0_0_in = 32'd0;
        A_sh_read0_0_write_en = 1'd0;
        A_sh_read0_0_clk = 1'd0;
        B0_0_addr0 = 4'd0;
        B0_0_addr1 = 4'd0;
        B0_0_write_data = 32'd0;
        B0_0_write_en = 1'd0;
        B0_0_clk = 1'd0;
        B_int_read0_0_in = 32'd0;
        B_int_read0_0_write_en = 1'd0;
        B_int_read0_0_clk = 1'd0;
        B_read0_0_in = 32'd0;
        B_read0_0_write_en = 1'd0;
        B_read0_0_clk = 1'd0;
        B_sh_read0_0_in = 32'd0;
        B_sh_read0_0_write_en = 1'd0;
        B_sh_read0_0_clk = 1'd0;
        C0_0_addr0 = 4'd0;
        C0_0_addr1 = 4'd0;
        C0_0_write_data = 32'd0;
        C0_0_write_en = 1'd0;
        C0_0_clk = 1'd0;
        C_int_read0_0_in = 32'd0;
        C_int_read0_0_write_en = 1'd0;
        C_int_read0_0_clk = 1'd0;
        C_read0_0_in = 32'd0;
        C_read0_0_write_en = 1'd0;
        C_read0_0_clk = 1'd0;
        C_sh_read0_0_in = 32'd0;
        C_sh_read0_0_write_en = 1'd0;
        C_sh_read0_0_clk = 1'd0;
        D0_0_addr0 = 4'd0;
        D0_0_addr1 = 4'd0;
        D0_0_write_data = 32'd0;
        D0_0_write_en = 1'd0;
        D0_0_clk = 1'd0;
        D_int_read0_0_in = 32'd0;
        D_int_read0_0_write_en = 1'd0;
        D_int_read0_0_clk = 1'd0;
        D_sh_read0_0_in = 32'd0;
        D_sh_read0_0_write_en = 1'd0;
        D_sh_read0_0_clk = 1'd0;
        add0_left = 4'd0;
        add0_right = 4'd0;
        add2_left = 32'd0;
        add2_right = 32'd0;
        alpha_int_read0_0_in = 32'd0;
        alpha_int_read0_0_write_en = 1'd0;
        alpha_int_read0_0_clk = 1'd0;
        beta_int_read0_0_in = 32'd0;
        beta_int_read0_0_write_en = 1'd0;
        beta_int_read0_0_clk = 1'd0;
        bin_read0_0_in = 32'd0;
        bin_read0_0_write_en = 1'd0;
        bin_read0_0_clk = 1'd0;
        bin_read1_0_in = 32'd0;
        bin_read1_0_write_en = 1'd0;
        bin_read1_0_clk = 1'd0;
        bin_read2_0_in = 32'd0;
        bin_read2_0_write_en = 1'd0;
        bin_read2_0_clk = 1'd0;
        bin_read3_0_in = 32'd0;
        bin_read3_0_write_en = 1'd0;
        bin_read3_0_clk = 1'd0;
        d_tmp_0_in = 32'd0;
        d_tmp_0_write_en = 1'd0;
        d_tmp_0_clk = 1'd0;
        i0_in = 4'd0;
        i0_write_en = 1'd0;
        i0_clk = 1'd0;
        i00_in = 4'd0;
        i00_write_en = 1'd0;
        i00_clk = 1'd0;
        i01_in = 4'd0;
        i01_write_en = 1'd0;
        i01_clk = 1'd0;
        i10_in = 4'd0;
        i10_write_en = 1'd0;
        i10_clk = 1'd0;
        j0_in = 4'd0;
        j0_write_en = 1'd0;
        j0_clk = 1'd0;
        j00_in = 4'd0;
        j00_write_en = 1'd0;
        j00_clk = 1'd0;
        j01_in = 4'd0;
        j01_write_en = 1'd0;
        j01_clk = 1'd0;
        j10_in = 4'd0;
        j10_write_en = 1'd0;
        j10_clk = 1'd0;
        k0_in = 4'd0;
        k0_write_en = 1'd0;
        k0_clk = 1'd0;
        k10_in = 4'd0;
        k10_write_en = 1'd0;
        k10_clk = 1'd0;
        le0_left = 4'd0;
        le0_right = 4'd0;
        mult_pipe0_left = 32'd0;
        mult_pipe0_right = 32'd0;
        mult_pipe0_go = 1'd0;
        mult_pipe0_clk = 1'd0;
        mult_pipe1_left = 32'd0;
        mult_pipe1_right = 32'd0;
        mult_pipe1_go = 1'd0;
        mult_pipe1_clk = 1'd0;
        mult_pipe2_left = 32'd0;
        mult_pipe2_right = 32'd0;
        mult_pipe2_go = 1'd0;
        mult_pipe2_clk = 1'd0;
        mult_pipe3_left = 32'd0;
        mult_pipe3_right = 32'd0;
        mult_pipe3_go = 1'd0;
        mult_pipe3_clk = 1'd0;
        rsh0_left = 4'd0;
        rsh0_right = 4'd0;
        rsh1_left = 4'd0;
        rsh1_right = 4'd0;
        tmp0_0_addr0 = 4'd0;
        tmp0_0_addr1 = 4'd0;
        tmp0_0_write_data = 32'd0;
        tmp0_0_write_en = 1'd0;
        tmp0_0_clk = 1'd0;
        tmp_int_read0_0_in = 32'd0;
        tmp_int_read0_0_write_en = 1'd0;
        tmp_int_read0_0_clk = 1'd0;
        tmp_read0_0_in = 32'd0;
        tmp_read0_0_write_en = 1'd0;
        tmp_read0_0_clk = 1'd0;
        tmp_sh_read0_0_in = 32'd0;
        tmp_sh_read0_0_write_en = 1'd0;
        tmp_sh_read0_0_clk = 1'd0;
        v1_0_in = 32'd0;
        v1_0_write_en = 1'd0;
        v1_0_clk = 1'd0;
        v_0_in = 32'd0;
        v_0_write_en = 1'd0;
        v_0_clk = 1'd0;
        par_reset_in = 1'd0;
        par_reset_write_en = 1'd0;
        par_reset_clk = 1'd0;
        par_done_reg_in = 1'd0;
        par_done_reg_write_en = 1'd0;
        par_done_reg_clk = 1'd0;
        par_done_reg0_in = 1'd0;
        par_done_reg0_write_en = 1'd0;
        par_done_reg0_clk = 1'd0;
        par_reset0_in = 1'd0;
        par_reset0_write_en = 1'd0;
        par_reset0_clk = 1'd0;
        par_done_reg1_in = 1'd0;
        par_done_reg1_write_en = 1'd0;
        par_done_reg1_clk = 1'd0;
        par_done_reg2_in = 1'd0;
        par_done_reg2_write_en = 1'd0;
        par_done_reg2_clk = 1'd0;
        par_reset1_in = 1'd0;
        par_reset1_write_en = 1'd0;
        par_reset1_clk = 1'd0;
        par_done_reg3_in = 1'd0;
        par_done_reg3_write_en = 1'd0;
        par_done_reg3_clk = 1'd0;
        par_done_reg4_in = 1'd0;
        par_done_reg4_write_en = 1'd0;
        par_done_reg4_clk = 1'd0;
        par_reset2_in = 1'd0;
        par_reset2_write_en = 1'd0;
        par_reset2_clk = 1'd0;
        par_done_reg5_in = 1'd0;
        par_done_reg5_write_en = 1'd0;
        par_done_reg5_clk = 1'd0;
        par_done_reg6_in = 1'd0;
        par_done_reg6_write_en = 1'd0;
        par_done_reg6_clk = 1'd0;
        fsm_in = 32'd0;
        fsm_write_en = 1'd0;
        fsm_clk = 1'd0;
        cond_computed_in = 1'd0;
        cond_computed_write_en = 1'd0;
        cond_computed_clk = 1'd0;
        cond_stored_in = 1'd0;
        cond_stored_write_en = 1'd0;
        cond_stored_clk = 1'd0;
        done_reg_in = 1'd0;
        done_reg_write_en = 1'd0;
        done_reg_clk = 1'd0;
        fsm0_in = 32'd0;
        fsm0_write_en = 1'd0;
        fsm0_clk = 1'd0;
        cond_computed0_in = 1'd0;
        cond_computed0_write_en = 1'd0;
        cond_computed0_clk = 1'd0;
        cond_stored0_in = 1'd0;
        cond_stored0_write_en = 1'd0;
        cond_stored0_clk = 1'd0;
        done_reg0_in = 1'd0;
        done_reg0_write_en = 1'd0;
        done_reg0_clk = 1'd0;
        par_reset3_in = 1'd0;
        par_reset3_write_en = 1'd0;
        par_reset3_clk = 1'd0;
        par_done_reg7_in = 1'd0;
        par_done_reg7_write_en = 1'd0;
        par_done_reg7_clk = 1'd0;
        par_done_reg8_in = 1'd0;
        par_done_reg8_write_en = 1'd0;
        par_done_reg8_clk = 1'd0;
        par_done_reg9_in = 1'd0;
        par_done_reg9_write_en = 1'd0;
        par_done_reg9_clk = 1'd0;
        fsm1_in = 32'd0;
        fsm1_write_en = 1'd0;
        fsm1_clk = 1'd0;
        cond_computed1_in = 1'd0;
        cond_computed1_write_en = 1'd0;
        cond_computed1_clk = 1'd0;
        cond_stored1_in = 1'd0;
        cond_stored1_write_en = 1'd0;
        cond_stored1_clk = 1'd0;
        done_reg1_in = 1'd0;
        done_reg1_write_en = 1'd0;
        done_reg1_clk = 1'd0;
        fsm2_in = 32'd0;
        fsm2_write_en = 1'd0;
        fsm2_clk = 1'd0;
        cond_computed2_in = 1'd0;
        cond_computed2_write_en = 1'd0;
        cond_computed2_clk = 1'd0;
        cond_stored2_in = 1'd0;
        cond_stored2_write_en = 1'd0;
        cond_stored2_clk = 1'd0;
        done_reg2_in = 1'd0;
        done_reg2_write_en = 1'd0;
        done_reg2_clk = 1'd0;
        fsm3_in = 32'd0;
        fsm3_write_en = 1'd0;
        fsm3_clk = 1'd0;
        cond_computed3_in = 1'd0;
        cond_computed3_write_en = 1'd0;
        cond_computed3_clk = 1'd0;
        cond_stored3_in = 1'd0;
        cond_stored3_write_en = 1'd0;
        cond_stored3_clk = 1'd0;
        done_reg3_in = 1'd0;
        done_reg3_write_en = 1'd0;
        done_reg3_clk = 1'd0;
        par_reset4_in = 1'd0;
        par_reset4_write_en = 1'd0;
        par_reset4_clk = 1'd0;
        par_done_reg10_in = 1'd0;
        par_done_reg10_write_en = 1'd0;
        par_done_reg10_clk = 1'd0;
        par_done_reg11_in = 1'd0;
        par_done_reg11_write_en = 1'd0;
        par_done_reg11_clk = 1'd0;
        fsm4_in = 32'd0;
        fsm4_write_en = 1'd0;
        fsm4_clk = 1'd0;
        cond_computed4_in = 1'd0;
        cond_computed4_write_en = 1'd0;
        cond_computed4_clk = 1'd0;
        cond_stored4_in = 1'd0;
        cond_stored4_write_en = 1'd0;
        cond_stored4_clk = 1'd0;
        done_reg4_in = 1'd0;
        done_reg4_write_en = 1'd0;
        done_reg4_clk = 1'd0;
        fsm5_in = 32'd0;
        fsm5_write_en = 1'd0;
        fsm5_clk = 1'd0;
        cond_computed5_in = 1'd0;
        cond_computed5_write_en = 1'd0;
        cond_computed5_clk = 1'd0;
        cond_stored5_in = 1'd0;
        cond_stored5_write_en = 1'd0;
        cond_stored5_clk = 1'd0;
        done_reg5_in = 1'd0;
        done_reg5_write_en = 1'd0;
        done_reg5_clk = 1'd0;
        fsm6_in = 32'd0;
        fsm6_write_en = 1'd0;
        fsm6_clk = 1'd0;
        cond_computed6_in = 1'd0;
        cond_computed6_write_en = 1'd0;
        cond_computed6_clk = 1'd0;
        cond_stored6_in = 1'd0;
        cond_stored6_write_en = 1'd0;
        cond_stored6_clk = 1'd0;
        done_reg6_in = 1'd0;
        done_reg6_write_en = 1'd0;
        done_reg6_clk = 1'd0;
        par_reset5_in = 1'd0;
        par_reset5_write_en = 1'd0;
        par_reset5_clk = 1'd0;
        par_done_reg12_in = 1'd0;
        par_done_reg12_write_en = 1'd0;
        par_done_reg12_clk = 1'd0;
        par_done_reg13_in = 1'd0;
        par_done_reg13_write_en = 1'd0;
        par_done_reg13_clk = 1'd0;
        par_reset6_in = 1'd0;
        par_reset6_write_en = 1'd0;
        par_reset6_clk = 1'd0;
        par_done_reg14_in = 1'd0;
        par_done_reg14_write_en = 1'd0;
        par_done_reg14_clk = 1'd0;
        par_done_reg15_in = 1'd0;
        par_done_reg15_write_en = 1'd0;
        par_done_reg15_clk = 1'd0;
        par_reset7_in = 1'd0;
        par_reset7_write_en = 1'd0;
        par_reset7_clk = 1'd0;
        par_done_reg16_in = 1'd0;
        par_done_reg16_write_en = 1'd0;
        par_done_reg16_clk = 1'd0;
        par_done_reg17_in = 1'd0;
        par_done_reg17_write_en = 1'd0;
        par_done_reg17_clk = 1'd0;
        par_reset8_in = 1'd0;
        par_reset8_write_en = 1'd0;
        par_reset8_clk = 1'd0;
        par_done_reg18_in = 1'd0;
        par_done_reg18_write_en = 1'd0;
        par_done_reg18_clk = 1'd0;
        par_done_reg19_in = 1'd0;
        par_done_reg19_write_en = 1'd0;
        par_done_reg19_clk = 1'd0;
        fsm7_in = 32'd0;
        fsm7_write_en = 1'd0;
        fsm7_clk = 1'd0;
        cond_computed7_in = 1'd0;
        cond_computed7_write_en = 1'd0;
        cond_computed7_clk = 1'd0;
        cond_stored7_in = 1'd0;
        cond_stored7_write_en = 1'd0;
        cond_stored7_clk = 1'd0;
        done_reg7_in = 1'd0;
        done_reg7_write_en = 1'd0;
        done_reg7_clk = 1'd0;
        fsm8_in = 32'd0;
        fsm8_write_en = 1'd0;
        fsm8_clk = 1'd0;
        cond_computed8_in = 1'd0;
        cond_computed8_write_en = 1'd0;
        cond_computed8_clk = 1'd0;
        cond_stored8_in = 1'd0;
        cond_stored8_write_en = 1'd0;
        cond_stored8_clk = 1'd0;
        done_reg8_in = 1'd0;
        done_reg8_write_en = 1'd0;
        done_reg8_clk = 1'd0;
        fsm9_in = 32'd0;
        fsm9_write_en = 1'd0;
        fsm9_clk = 1'd0;
    end
    std_mem_d2 # (
        .d0_idx_size(4),
        .d0_size(8),
        .d1_idx_size(4),
        .d1_size(8),
        .width(32)
    ) A0_0 (
        .addr0(A0_0_addr0),
        .addr1(A0_0_addr1),
        .clk(A0_0_clk),
        .done(A0_0_done),
        .read_data(A0_0_read_data),
        .write_data(A0_0_write_data),
        .write_en(A0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_int_read0_0 (
        .clk(A_int_read0_0_clk),
        .done(A_int_read0_0_done),
        .in(A_int_read0_0_in),
        .out(A_int_read0_0_out),
        .write_en(A_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_read0_0 (
        .clk(A_read0_0_clk),
        .done(A_read0_0_done),
        .in(A_read0_0_in),
        .out(A_read0_0_out),
        .write_en(A_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) A_sh_read0_0 (
        .clk(A_sh_read0_0_clk),
        .done(A_sh_read0_0_done),
        .in(A_sh_read0_0_in),
        .out(A_sh_read0_0_out),
        .write_en(A_sh_read0_0_write_en)
    );
    std_mem_d2 # (
        .d0_idx_size(4),
        .d0_size(8),
        .d1_idx_size(4),
        .d1_size(8),
        .width(32)
    ) B0_0 (
        .addr0(B0_0_addr0),
        .addr1(B0_0_addr1),
        .clk(B0_0_clk),
        .done(B0_0_done),
        .read_data(B0_0_read_data),
        .write_data(B0_0_write_data),
        .write_en(B0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) B_int_read0_0 (
        .clk(B_int_read0_0_clk),
        .done(B_int_read0_0_done),
        .in(B_int_read0_0_in),
        .out(B_int_read0_0_out),
        .write_en(B_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) B_read0_0 (
        .clk(B_read0_0_clk),
        .done(B_read0_0_done),
        .in(B_read0_0_in),
        .out(B_read0_0_out),
        .write_en(B_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) B_sh_read0_0 (
        .clk(B_sh_read0_0_clk),
        .done(B_sh_read0_0_done),
        .in(B_sh_read0_0_in),
        .out(B_sh_read0_0_out),
        .write_en(B_sh_read0_0_write_en)
    );
    std_mem_d2 # (
        .d0_idx_size(4),
        .d0_size(8),
        .d1_idx_size(4),
        .d1_size(8),
        .width(32)
    ) C0_0 (
        .addr0(C0_0_addr0),
        .addr1(C0_0_addr1),
        .clk(C0_0_clk),
        .done(C0_0_done),
        .read_data(C0_0_read_data),
        .write_data(C0_0_write_data),
        .write_en(C0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) C_int_read0_0 (
        .clk(C_int_read0_0_clk),
        .done(C_int_read0_0_done),
        .in(C_int_read0_0_in),
        .out(C_int_read0_0_out),
        .write_en(C_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) C_read0_0 (
        .clk(C_read0_0_clk),
        .done(C_read0_0_done),
        .in(C_read0_0_in),
        .out(C_read0_0_out),
        .write_en(C_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) C_sh_read0_0 (
        .clk(C_sh_read0_0_clk),
        .done(C_sh_read0_0_done),
        .in(C_sh_read0_0_in),
        .out(C_sh_read0_0_out),
        .write_en(C_sh_read0_0_write_en)
    );
    std_mem_d2 # (
        .d0_idx_size(4),
        .d0_size(8),
        .d1_idx_size(4),
        .d1_size(8),
        .width(32)
    ) D0_0 (
        .addr0(D0_0_addr0),
        .addr1(D0_0_addr1),
        .clk(D0_0_clk),
        .done(D0_0_done),
        .read_data(D0_0_read_data),
        .write_data(D0_0_write_data),
        .write_en(D0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) D_int_read0_0 (
        .clk(D_int_read0_0_clk),
        .done(D_int_read0_0_done),
        .in(D_int_read0_0_in),
        .out(D_int_read0_0_out),
        .write_en(D_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) D_sh_read0_0 (
        .clk(D_sh_read0_0_clk),
        .done(D_sh_read0_0_done),
        .in(D_sh_read0_0_in),
        .out(D_sh_read0_0_out),
        .write_en(D_sh_read0_0_write_en)
    );
    std_add # (
        .width(4)
    ) add0 (
        .left(add0_left),
        .out(add0_out),
        .right(add0_right)
    );
    std_add # (
        .width(32)
    ) add2 (
        .left(add2_left),
        .out(add2_out),
        .right(add2_right)
    );
    std_reg # (
        .width(32)
    ) alpha_int_read0_0 (
        .clk(alpha_int_read0_0_clk),
        .done(alpha_int_read0_0_done),
        .in(alpha_int_read0_0_in),
        .out(alpha_int_read0_0_out),
        .write_en(alpha_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) beta_int_read0_0 (
        .clk(beta_int_read0_0_clk),
        .done(beta_int_read0_0_done),
        .in(beta_int_read0_0_in),
        .out(beta_int_read0_0_out),
        .write_en(beta_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read0_0 (
        .clk(bin_read0_0_clk),
        .done(bin_read0_0_done),
        .in(bin_read0_0_in),
        .out(bin_read0_0_out),
        .write_en(bin_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read1_0 (
        .clk(bin_read1_0_clk),
        .done(bin_read1_0_done),
        .in(bin_read1_0_in),
        .out(bin_read1_0_out),
        .write_en(bin_read1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read2_0 (
        .clk(bin_read2_0_clk),
        .done(bin_read2_0_done),
        .in(bin_read2_0_in),
        .out(bin_read2_0_out),
        .write_en(bin_read2_0_write_en)
    );
    std_reg # (
        .width(32)
    ) bin_read3_0 (
        .clk(bin_read3_0_clk),
        .done(bin_read3_0_done),
        .in(bin_read3_0_in),
        .out(bin_read3_0_out),
        .write_en(bin_read3_0_write_en)
    );
    std_const # (
        .value(0),
        .width(4)
    ) const0 (
        .out(const0_out)
    );
    std_const # (
        .value(7),
        .width(4)
    ) const1 (
        .out(const1_out)
    );
    std_const # (
        .value(0),
        .width(4)
    ) const10 (
        .out(const10_out)
    );
    std_const # (
        .value(1),
        .width(4)
    ) const14 (
        .out(const14_out)
    );
    std_const # (
        .value(0),
        .width(32)
    ) const20 (
        .out(const20_out)
    );
    std_const # (
        .value(0),
        .width(1)
    ) const23 (
        .out(const23_out)
    );
    std_reg # (
        .width(32)
    ) d_tmp_0 (
        .clk(d_tmp_0_clk),
        .done(d_tmp_0_done),
        .in(d_tmp_0_in),
        .out(d_tmp_0_out),
        .write_en(d_tmp_0_write_en)
    );
    std_reg # (
        .width(4)
    ) i0 (
        .clk(i0_clk),
        .done(i0_done),
        .in(i0_in),
        .out(i0_out),
        .write_en(i0_write_en)
    );
    std_reg # (
        .width(4)
    ) i00 (
        .clk(i00_clk),
        .done(i00_done),
        .in(i00_in),
        .out(i00_out),
        .write_en(i00_write_en)
    );
    std_reg # (
        .width(4)
    ) i01 (
        .clk(i01_clk),
        .done(i01_done),
        .in(i01_in),
        .out(i01_out),
        .write_en(i01_write_en)
    );
    std_reg # (
        .width(4)
    ) i10 (
        .clk(i10_clk),
        .done(i10_done),
        .in(i10_in),
        .out(i10_out),
        .write_en(i10_write_en)
    );
    std_reg # (
        .width(4)
    ) j0 (
        .clk(j0_clk),
        .done(j0_done),
        .in(j0_in),
        .out(j0_out),
        .write_en(j0_write_en)
    );
    std_reg # (
        .width(4)
    ) j00 (
        .clk(j00_clk),
        .done(j00_done),
        .in(j00_in),
        .out(j00_out),
        .write_en(j00_write_en)
    );
    std_reg # (
        .width(4)
    ) j01 (
        .clk(j01_clk),
        .done(j01_done),
        .in(j01_in),
        .out(j01_out),
        .write_en(j01_write_en)
    );
    std_reg # (
        .width(4)
    ) j10 (
        .clk(j10_clk),
        .done(j10_done),
        .in(j10_in),
        .out(j10_out),
        .write_en(j10_write_en)
    );
    std_reg # (
        .width(4)
    ) k0 (
        .clk(k0_clk),
        .done(k0_done),
        .in(k0_in),
        .out(k0_out),
        .write_en(k0_write_en)
    );
    std_reg # (
        .width(4)
    ) k10 (
        .clk(k10_clk),
        .done(k10_done),
        .in(k10_in),
        .out(k10_out),
        .write_en(k10_write_en)
    );
    std_le # (
        .width(4)
    ) le0 (
        .left(le0_left),
        .out(le0_out),
        .right(le0_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe0 (
        .clk(mult_pipe0_clk),
        .done(mult_pipe0_done),
        .go(mult_pipe0_go),
        .left(mult_pipe0_left),
        .out(mult_pipe0_out),
        .right(mult_pipe0_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe1 (
        .clk(mult_pipe1_clk),
        .done(mult_pipe1_done),
        .go(mult_pipe1_go),
        .left(mult_pipe1_left),
        .out(mult_pipe1_out),
        .right(mult_pipe1_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe2 (
        .clk(mult_pipe2_clk),
        .done(mult_pipe2_done),
        .go(mult_pipe2_go),
        .left(mult_pipe2_left),
        .out(mult_pipe2_out),
        .right(mult_pipe2_right)
    );
    std_mult_pipe # (
        .width(32)
    ) mult_pipe3 (
        .clk(mult_pipe3_clk),
        .done(mult_pipe3_done),
        .go(mult_pipe3_go),
        .left(mult_pipe3_left),
        .out(mult_pipe3_out),
        .right(mult_pipe3_right)
    );
    std_rsh # (
        .width(4)
    ) rsh0 (
        .left(rsh0_left),
        .out(rsh0_out),
        .right(rsh0_right)
    );
    std_rsh # (
        .width(4)
    ) rsh1 (
        .left(rsh1_left),
        .out(rsh1_out),
        .right(rsh1_right)
    );
    std_mem_d2 # (
        .d0_idx_size(4),
        .d0_size(8),
        .d1_idx_size(4),
        .d1_size(8),
        .width(32)
    ) tmp0_0 (
        .addr0(tmp0_0_addr0),
        .addr1(tmp0_0_addr1),
        .clk(tmp0_0_clk),
        .done(tmp0_0_done),
        .read_data(tmp0_0_read_data),
        .write_data(tmp0_0_write_data),
        .write_en(tmp0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) tmp_int_read0_0 (
        .clk(tmp_int_read0_0_clk),
        .done(tmp_int_read0_0_done),
        .in(tmp_int_read0_0_in),
        .out(tmp_int_read0_0_out),
        .write_en(tmp_int_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) tmp_read0_0 (
        .clk(tmp_read0_0_clk),
        .done(tmp_read0_0_done),
        .in(tmp_read0_0_in),
        .out(tmp_read0_0_out),
        .write_en(tmp_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) tmp_sh_read0_0 (
        .clk(tmp_sh_read0_0_clk),
        .done(tmp_sh_read0_0_done),
        .in(tmp_sh_read0_0_in),
        .out(tmp_sh_read0_0_out),
        .write_en(tmp_sh_read0_0_write_en)
    );
    std_reg # (
        .width(32)
    ) v1_0 (
        .clk(v1_0_clk),
        .done(v1_0_done),
        .in(v1_0_in),
        .out(v1_0_out),
        .write_en(v1_0_write_en)
    );
    std_reg # (
        .width(32)
    ) v_0 (
        .clk(v_0_clk),
        .done(v_0_done),
        .in(v_0_in),
        .out(v_0_out),
        .write_en(v_0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset (
        .clk(par_reset_clk),
        .done(par_reset_done),
        .in(par_reset_in),
        .out(par_reset_out),
        .write_en(par_reset_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg (
        .clk(par_done_reg_clk),
        .done(par_done_reg_done),
        .in(par_done_reg_in),
        .out(par_done_reg_out),
        .write_en(par_done_reg_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg0 (
        .clk(par_done_reg0_clk),
        .done(par_done_reg0_done),
        .in(par_done_reg0_in),
        .out(par_done_reg0_out),
        .write_en(par_done_reg0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset0 (
        .clk(par_reset0_clk),
        .done(par_reset0_done),
        .in(par_reset0_in),
        .out(par_reset0_out),
        .write_en(par_reset0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg1 (
        .clk(par_done_reg1_clk),
        .done(par_done_reg1_done),
        .in(par_done_reg1_in),
        .out(par_done_reg1_out),
        .write_en(par_done_reg1_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg2 (
        .clk(par_done_reg2_clk),
        .done(par_done_reg2_done),
        .in(par_done_reg2_in),
        .out(par_done_reg2_out),
        .write_en(par_done_reg2_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset1 (
        .clk(par_reset1_clk),
        .done(par_reset1_done),
        .in(par_reset1_in),
        .out(par_reset1_out),
        .write_en(par_reset1_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg3 (
        .clk(par_done_reg3_clk),
        .done(par_done_reg3_done),
        .in(par_done_reg3_in),
        .out(par_done_reg3_out),
        .write_en(par_done_reg3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg4 (
        .clk(par_done_reg4_clk),
        .done(par_done_reg4_done),
        .in(par_done_reg4_in),
        .out(par_done_reg4_out),
        .write_en(par_done_reg4_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset2 (
        .clk(par_reset2_clk),
        .done(par_reset2_done),
        .in(par_reset2_in),
        .out(par_reset2_out),
        .write_en(par_reset2_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg5 (
        .clk(par_done_reg5_clk),
        .done(par_done_reg5_done),
        .in(par_done_reg5_in),
        .out(par_done_reg5_out),
        .write_en(par_done_reg5_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg6 (
        .clk(par_done_reg6_clk),
        .done(par_done_reg6_done),
        .in(par_done_reg6_in),
        .out(par_done_reg6_out),
        .write_en(par_done_reg6_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm (
        .clk(fsm_clk),
        .done(fsm_done),
        .in(fsm_in),
        .out(fsm_out),
        .write_en(fsm_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed (
        .clk(cond_computed_clk),
        .done(cond_computed_done),
        .in(cond_computed_in),
        .out(cond_computed_out),
        .write_en(cond_computed_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored (
        .clk(cond_stored_clk),
        .done(cond_stored_done),
        .in(cond_stored_in),
        .out(cond_stored_out),
        .write_en(cond_stored_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg (
        .clk(done_reg_clk),
        .done(done_reg_done),
        .in(done_reg_in),
        .out(done_reg_out),
        .write_en(done_reg_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm0 (
        .clk(fsm0_clk),
        .done(fsm0_done),
        .in(fsm0_in),
        .out(fsm0_out),
        .write_en(fsm0_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed0 (
        .clk(cond_computed0_clk),
        .done(cond_computed0_done),
        .in(cond_computed0_in),
        .out(cond_computed0_out),
        .write_en(cond_computed0_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored0 (
        .clk(cond_stored0_clk),
        .done(cond_stored0_done),
        .in(cond_stored0_in),
        .out(cond_stored0_out),
        .write_en(cond_stored0_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg0 (
        .clk(done_reg0_clk),
        .done(done_reg0_done),
        .in(done_reg0_in),
        .out(done_reg0_out),
        .write_en(done_reg0_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset3 (
        .clk(par_reset3_clk),
        .done(par_reset3_done),
        .in(par_reset3_in),
        .out(par_reset3_out),
        .write_en(par_reset3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg7 (
        .clk(par_done_reg7_clk),
        .done(par_done_reg7_done),
        .in(par_done_reg7_in),
        .out(par_done_reg7_out),
        .write_en(par_done_reg7_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg8 (
        .clk(par_done_reg8_clk),
        .done(par_done_reg8_done),
        .in(par_done_reg8_in),
        .out(par_done_reg8_out),
        .write_en(par_done_reg8_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg9 (
        .clk(par_done_reg9_clk),
        .done(par_done_reg9_done),
        .in(par_done_reg9_in),
        .out(par_done_reg9_out),
        .write_en(par_done_reg9_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm1 (
        .clk(fsm1_clk),
        .done(fsm1_done),
        .in(fsm1_in),
        .out(fsm1_out),
        .write_en(fsm1_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed1 (
        .clk(cond_computed1_clk),
        .done(cond_computed1_done),
        .in(cond_computed1_in),
        .out(cond_computed1_out),
        .write_en(cond_computed1_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored1 (
        .clk(cond_stored1_clk),
        .done(cond_stored1_done),
        .in(cond_stored1_in),
        .out(cond_stored1_out),
        .write_en(cond_stored1_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg1 (
        .clk(done_reg1_clk),
        .done(done_reg1_done),
        .in(done_reg1_in),
        .out(done_reg1_out),
        .write_en(done_reg1_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm2 (
        .clk(fsm2_clk),
        .done(fsm2_done),
        .in(fsm2_in),
        .out(fsm2_out),
        .write_en(fsm2_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed2 (
        .clk(cond_computed2_clk),
        .done(cond_computed2_done),
        .in(cond_computed2_in),
        .out(cond_computed2_out),
        .write_en(cond_computed2_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored2 (
        .clk(cond_stored2_clk),
        .done(cond_stored2_done),
        .in(cond_stored2_in),
        .out(cond_stored2_out),
        .write_en(cond_stored2_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg2 (
        .clk(done_reg2_clk),
        .done(done_reg2_done),
        .in(done_reg2_in),
        .out(done_reg2_out),
        .write_en(done_reg2_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm3 (
        .clk(fsm3_clk),
        .done(fsm3_done),
        .in(fsm3_in),
        .out(fsm3_out),
        .write_en(fsm3_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed3 (
        .clk(cond_computed3_clk),
        .done(cond_computed3_done),
        .in(cond_computed3_in),
        .out(cond_computed3_out),
        .write_en(cond_computed3_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored3 (
        .clk(cond_stored3_clk),
        .done(cond_stored3_done),
        .in(cond_stored3_in),
        .out(cond_stored3_out),
        .write_en(cond_stored3_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg3 (
        .clk(done_reg3_clk),
        .done(done_reg3_done),
        .in(done_reg3_in),
        .out(done_reg3_out),
        .write_en(done_reg3_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset4 (
        .clk(par_reset4_clk),
        .done(par_reset4_done),
        .in(par_reset4_in),
        .out(par_reset4_out),
        .write_en(par_reset4_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg10 (
        .clk(par_done_reg10_clk),
        .done(par_done_reg10_done),
        .in(par_done_reg10_in),
        .out(par_done_reg10_out),
        .write_en(par_done_reg10_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg11 (
        .clk(par_done_reg11_clk),
        .done(par_done_reg11_done),
        .in(par_done_reg11_in),
        .out(par_done_reg11_out),
        .write_en(par_done_reg11_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm4 (
        .clk(fsm4_clk),
        .done(fsm4_done),
        .in(fsm4_in),
        .out(fsm4_out),
        .write_en(fsm4_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed4 (
        .clk(cond_computed4_clk),
        .done(cond_computed4_done),
        .in(cond_computed4_in),
        .out(cond_computed4_out),
        .write_en(cond_computed4_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored4 (
        .clk(cond_stored4_clk),
        .done(cond_stored4_done),
        .in(cond_stored4_in),
        .out(cond_stored4_out),
        .write_en(cond_stored4_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg4 (
        .clk(done_reg4_clk),
        .done(done_reg4_done),
        .in(done_reg4_in),
        .out(done_reg4_out),
        .write_en(done_reg4_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm5 (
        .clk(fsm5_clk),
        .done(fsm5_done),
        .in(fsm5_in),
        .out(fsm5_out),
        .write_en(fsm5_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed5 (
        .clk(cond_computed5_clk),
        .done(cond_computed5_done),
        .in(cond_computed5_in),
        .out(cond_computed5_out),
        .write_en(cond_computed5_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored5 (
        .clk(cond_stored5_clk),
        .done(cond_stored5_done),
        .in(cond_stored5_in),
        .out(cond_stored5_out),
        .write_en(cond_stored5_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg5 (
        .clk(done_reg5_clk),
        .done(done_reg5_done),
        .in(done_reg5_in),
        .out(done_reg5_out),
        .write_en(done_reg5_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm6 (
        .clk(fsm6_clk),
        .done(fsm6_done),
        .in(fsm6_in),
        .out(fsm6_out),
        .write_en(fsm6_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed6 (
        .clk(cond_computed6_clk),
        .done(cond_computed6_done),
        .in(cond_computed6_in),
        .out(cond_computed6_out),
        .write_en(cond_computed6_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored6 (
        .clk(cond_stored6_clk),
        .done(cond_stored6_done),
        .in(cond_stored6_in),
        .out(cond_stored6_out),
        .write_en(cond_stored6_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg6 (
        .clk(done_reg6_clk),
        .done(done_reg6_done),
        .in(done_reg6_in),
        .out(done_reg6_out),
        .write_en(done_reg6_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset5 (
        .clk(par_reset5_clk),
        .done(par_reset5_done),
        .in(par_reset5_in),
        .out(par_reset5_out),
        .write_en(par_reset5_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg12 (
        .clk(par_done_reg12_clk),
        .done(par_done_reg12_done),
        .in(par_done_reg12_in),
        .out(par_done_reg12_out),
        .write_en(par_done_reg12_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg13 (
        .clk(par_done_reg13_clk),
        .done(par_done_reg13_done),
        .in(par_done_reg13_in),
        .out(par_done_reg13_out),
        .write_en(par_done_reg13_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset6 (
        .clk(par_reset6_clk),
        .done(par_reset6_done),
        .in(par_reset6_in),
        .out(par_reset6_out),
        .write_en(par_reset6_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg14 (
        .clk(par_done_reg14_clk),
        .done(par_done_reg14_done),
        .in(par_done_reg14_in),
        .out(par_done_reg14_out),
        .write_en(par_done_reg14_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg15 (
        .clk(par_done_reg15_clk),
        .done(par_done_reg15_done),
        .in(par_done_reg15_in),
        .out(par_done_reg15_out),
        .write_en(par_done_reg15_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset7 (
        .clk(par_reset7_clk),
        .done(par_reset7_done),
        .in(par_reset7_in),
        .out(par_reset7_out),
        .write_en(par_reset7_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg16 (
        .clk(par_done_reg16_clk),
        .done(par_done_reg16_done),
        .in(par_done_reg16_in),
        .out(par_done_reg16_out),
        .write_en(par_done_reg16_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg17 (
        .clk(par_done_reg17_clk),
        .done(par_done_reg17_done),
        .in(par_done_reg17_in),
        .out(par_done_reg17_out),
        .write_en(par_done_reg17_write_en)
    );
    std_reg # (
        .width(1)
    ) par_reset8 (
        .clk(par_reset8_clk),
        .done(par_reset8_done),
        .in(par_reset8_in),
        .out(par_reset8_out),
        .write_en(par_reset8_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg18 (
        .clk(par_done_reg18_clk),
        .done(par_done_reg18_done),
        .in(par_done_reg18_in),
        .out(par_done_reg18_out),
        .write_en(par_done_reg18_write_en)
    );
    std_reg # (
        .width(1)
    ) par_done_reg19 (
        .clk(par_done_reg19_clk),
        .done(par_done_reg19_done),
        .in(par_done_reg19_in),
        .out(par_done_reg19_out),
        .write_en(par_done_reg19_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm7 (
        .clk(fsm7_clk),
        .done(fsm7_done),
        .in(fsm7_in),
        .out(fsm7_out),
        .write_en(fsm7_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed7 (
        .clk(cond_computed7_clk),
        .done(cond_computed7_done),
        .in(cond_computed7_in),
        .out(cond_computed7_out),
        .write_en(cond_computed7_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored7 (
        .clk(cond_stored7_clk),
        .done(cond_stored7_done),
        .in(cond_stored7_in),
        .out(cond_stored7_out),
        .write_en(cond_stored7_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg7 (
        .clk(done_reg7_clk),
        .done(done_reg7_done),
        .in(done_reg7_in),
        .out(done_reg7_out),
        .write_en(done_reg7_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm8 (
        .clk(fsm8_clk),
        .done(fsm8_done),
        .in(fsm8_in),
        .out(fsm8_out),
        .write_en(fsm8_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_computed8 (
        .clk(cond_computed8_clk),
        .done(cond_computed8_done),
        .in(cond_computed8_in),
        .out(cond_computed8_out),
        .write_en(cond_computed8_write_en)
    );
    std_reg # (
        .width(1)
    ) cond_stored8 (
        .clk(cond_stored8_clk),
        .done(cond_stored8_done),
        .in(cond_stored8_in),
        .out(cond_stored8_out),
        .write_en(cond_stored8_write_en)
    );
    std_reg # (
        .width(1)
    ) done_reg8 (
        .clk(done_reg8_clk),
        .done(done_reg8_done),
        .in(done_reg8_in),
        .out(done_reg8_out),
        .write_en(done_reg8_write_en)
    );
    std_reg # (
        .width(32)
    ) fsm9 (
        .clk(fsm9_clk),
        .done(fsm9_done),
        .in(fsm9_in),
        .out(fsm9_out),
        .write_en(fsm9_write_en)
    );
    always_comb begin
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            A0_0_addr0 = rsh1_out;
        end else if((~(par_done_reg8_out | A_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            A0_0_addr0 = i0_out;
        end else if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            A0_0_addr0 = rsh1_out;
        end else A0_0_addr0 = 4'd0;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            A0_0_addr1 = rsh0_out;
        end else if((~(par_done_reg8_out | A_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            A0_0_addr1 = k0_out;
        end else if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            A0_0_addr1 = rsh0_out;
        end else A0_0_addr1 = 4'd0;
        A0_0_clk = clk;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            A0_0_write_data = A_int_read0_0_out;
        end else A0_0_write_data = 32'd0;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            A0_0_write_en = 1'd1;
        end else A0_0_write_en = 1'd0;
        A_int_read0_0_clk = clk;
        if((((fsm_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            A_int_read0_0_in = A_int0_0_read_data;
        end else A_int_read0_0_in = 32'd0;
        if((((fsm_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            A_int_read0_0_write_en = 1'd1;
        end else A_int_read0_0_write_en = 1'd0;
        A_read0_0_clk = clk;
        if((~(par_done_reg8_out | A_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            A_read0_0_in = A0_0_read_data;
        end else A_read0_0_in = 32'd0;
        if((~(par_done_reg8_out | A_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            A_read0_0_write_en = 1'd1;
        end else A_read0_0_write_en = 1'd0;
        A_sh_read0_0_clk = clk;
        if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            A_sh_read0_0_in = A0_0_read_data;
        end else A_sh_read0_0_in = 32'd0;
        if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            A_sh_read0_0_write_en = 1'd1;
        end else A_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg9_out | B_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            B0_0_addr0 = k0_out;
        end else if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B0_0_addr0 = rsh1_out;
        end else if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B0_0_addr0 = rsh1_out;
        end else B0_0_addr0 = 4'd0;
        if((~(par_done_reg9_out | B_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            B0_0_addr1 = j0_out;
        end else if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B0_0_addr1 = rsh0_out;
        end else if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B0_0_addr1 = rsh0_out;
        end else B0_0_addr1 = 4'd0;
        B0_0_clk = clk;
        if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B0_0_write_data = B_int_read0_0_out;
        end else B0_0_write_data = 32'd0;
        if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B0_0_write_en = 1'd1;
        end else B0_0_write_en = 1'd0;
        B_int_read0_0_clk = clk;
        if((~(par_done_reg0_out | B_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B_int_read0_0_in = B_int0_0_read_data;
        end else B_int_read0_0_in = 32'd0;
        if((~(par_done_reg0_out | B_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B_int_read0_0_write_en = 1'd1;
        end else B_int_read0_0_write_en = 1'd0;
        B_read0_0_clk = clk;
        if((~(par_done_reg9_out | B_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            B_read0_0_in = B0_0_read_data;
        end else B_read0_0_in = 32'd0;
        if((~(par_done_reg9_out | B_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            B_read0_0_write_en = 1'd1;
        end else B_read0_0_write_en = 1'd0;
        B_sh_read0_0_clk = clk;
        if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B_sh_read0_0_in = B0_0_read_data;
        end else B_sh_read0_0_in = 32'd0;
        if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B_sh_read0_0_write_en = 1'd1;
        end else B_sh_read0_0_write_en = 1'd0;
        if((~(par_done_reg11_out | C_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            C0_0_addr0 = k10_out;
        end else if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C0_0_addr0 = rsh1_out;
        end else if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C0_0_addr0 = rsh1_out;
        end else C0_0_addr0 = 4'd0;
        if((~(par_done_reg11_out | C_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            C0_0_addr1 = j10_out;
        end else if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C0_0_addr1 = rsh0_out;
        end else if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C0_0_addr1 = rsh0_out;
        end else C0_0_addr1 = 4'd0;
        C0_0_clk = clk;
        if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C0_0_write_data = C_int_read0_0_out;
        end else C0_0_write_data = 32'd0;
        if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C0_0_write_en = 1'd1;
        end else C0_0_write_en = 1'd0;
        C_int_read0_0_clk = clk;
        if((~(par_done_reg2_out | C_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C_int_read0_0_in = C_int0_0_read_data;
        end else C_int_read0_0_in = 32'd0;
        if((~(par_done_reg2_out | C_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C_int_read0_0_write_en = 1'd1;
        end else C_int_read0_0_write_en = 1'd0;
        C_read0_0_clk = clk;
        if((~(par_done_reg11_out | C_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            C_read0_0_in = C0_0_read_data;
        end else C_read0_0_in = 32'd0;
        if((~(par_done_reg11_out | C_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            C_read0_0_write_en = 1'd1;
        end else C_read0_0_write_en = 1'd0;
        C_sh_read0_0_clk = clk;
        if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C_sh_read0_0_in = C0_0_read_data;
        end else C_sh_read0_0_in = 32'd0;
        if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C_sh_read0_0_write_en = 1'd1;
        end else C_sh_read0_0_write_en = 1'd0;
        if((((fsm5_out == 32'd0) & ~d_tmp_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            D0_0_addr0 = i10_out;
        end else if((((fsm5_out == 32'd3) & ~D0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            D0_0_addr0 = i10_out;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            D0_0_addr0 = i10_out;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            D0_0_addr0 = i10_out;
        end else if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D0_0_addr0 = rsh1_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D0_0_addr0 = rsh1_out;
        end else D0_0_addr0 = 4'd0;
        if((((fsm5_out == 32'd0) & ~d_tmp_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            D0_0_addr1 = j10_out;
        end else if((((fsm5_out == 32'd3) & ~D0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            D0_0_addr1 = j10_out;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            D0_0_addr1 = j10_out;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            D0_0_addr1 = j10_out;
        end else if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D0_0_addr1 = rsh0_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D0_0_addr1 = rsh0_out;
        end else D0_0_addr1 = 4'd0;
        D0_0_clk = clk;
        if((((fsm5_out == 32'd3) & ~D0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            D0_0_write_data = bin_read2_0_out;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            D0_0_write_data = add2_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D0_0_write_data = D_int_read0_0_out;
        end else D0_0_write_data = 32'd0;
        if((((fsm5_out == 32'd3) & ~D0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            D0_0_write_en = 1'd1;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            D0_0_write_en = 1'd1;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D0_0_write_en = 1'd1;
        end else D0_0_write_en = 1'd0;
        D_int_read0_0_clk = clk;
        if((~(par_done_reg4_out | D_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D_int_read0_0_in = D_int0_0_read_data;
        end else D_int_read0_0_in = 32'd0;
        if((~(par_done_reg4_out | D_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D_int_read0_0_write_en = 1'd1;
        end else D_int_read0_0_write_en = 1'd0;
        D_sh_read0_0_clk = clk;
        if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D_sh_read0_0_in = D0_0_read_data;
        end else D_sh_read0_0_in = 32'd0;
        if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D_sh_read0_0_write_en = 1'd1;
        end else D_sh_read0_0_write_en = 1'd0;
        if((((fsm_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            A_int0_0_addr0 = i00_out;
        end else if((~(par_done_reg12_out | A_int0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            A_int0_0_addr0 = i01_out;
        end else A_int0_0_addr0 = 4'd0;
        if((((fsm_out == 32'd0) & ~A_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            A_int0_0_addr1 = j00_out;
        end else if((~(par_done_reg12_out | A_int0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            A_int0_0_addr1 = j01_out;
        end else A_int0_0_addr1 = 4'd0;
        A_int0_0_clk = clk;
        if((~(par_done_reg12_out | A_int0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            A_int0_0_write_data = A_sh_read0_0_out;
        end else A_int0_0_write_data = 32'd0;
        if((~(par_done_reg12_out | A_int0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            A_int0_0_write_en = 1'd1;
        end else A_int0_0_write_en = 1'd0;
        if((~(par_done_reg0_out | B_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B_int0_0_addr0 = i00_out;
        end else if((~(par_done_reg14_out | B_int0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B_int0_0_addr0 = i01_out;
        end else B_int0_0_addr0 = 4'd0;
        if((~(par_done_reg0_out | B_int_read0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            B_int0_0_addr1 = j00_out;
        end else if((~(par_done_reg14_out | B_int0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B_int0_0_addr1 = j01_out;
        end else B_int0_0_addr1 = 4'd0;
        B_int0_0_clk = clk;
        if((~(par_done_reg14_out | B_int0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B_int0_0_write_data = B_sh_read0_0_out;
        end else B_int0_0_write_data = 32'd0;
        if((~(par_done_reg14_out | B_int0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            B_int0_0_write_en = 1'd1;
        end else B_int0_0_write_en = 1'd0;
        if((~(par_done_reg16_out | C_int0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C_int0_0_addr0 = i01_out;
        end else if((~(par_done_reg2_out | C_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C_int0_0_addr0 = i00_out;
        end else C_int0_0_addr0 = 4'd0;
        if((~(par_done_reg16_out | C_int0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C_int0_0_addr1 = j01_out;
        end else if((~(par_done_reg2_out | C_int_read0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            C_int0_0_addr1 = j00_out;
        end else C_int0_0_addr1 = 4'd0;
        C_int0_0_clk = clk;
        if((~(par_done_reg16_out | C_int0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C_int0_0_write_data = C_sh_read0_0_out;
        end else C_int0_0_write_data = 32'd0;
        if((~(par_done_reg16_out | C_int0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            C_int0_0_write_en = 1'd1;
        end else C_int0_0_write_en = 1'd0;
        if((~(par_done_reg18_out | D_int0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D_int0_0_addr0 = i01_out;
        end else if((~(par_done_reg4_out | D_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D_int0_0_addr0 = i00_out;
        end else D_int0_0_addr0 = 4'd0;
        if((~(par_done_reg18_out | D_int0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D_int0_0_addr1 = j01_out;
        end else if((~(par_done_reg4_out | D_int_read0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            D_int0_0_addr1 = j00_out;
        end else D_int0_0_addr1 = 4'd0;
        D_int0_0_clk = clk;
        if((~(par_done_reg18_out | D_int0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D_int0_0_write_data = D_sh_read0_0_out;
        end else D_int0_0_write_data = 32'd0;
        if((~(par_done_reg18_out | D_int0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            D_int0_0_write_en = 1'd1;
        end else D_int0_0_write_en = 1'd0;
        if((~(par_done_reg7_out | alpha_int_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            alpha_int0_addr0 = const23_out;
        end else alpha_int0_addr0 = 1'd0;
        alpha_int0_clk = clk;
        if((((fsm5_out == 32'd1) & ~beta_int_read0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            beta_int0_addr0 = const23_out;
        end else beta_int0_addr0 = 1'd0;
        beta_int0_clk = clk;
        if((fsm9_out == 32'd8)) begin
            done = 1'd1;
        end else if((fsm9_out == 32'd8)) begin
            done = 1'd1;
        end else done = 1'd0;
        if((((fsm7_out == 32'd5) & ~tmp_int0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            tmp_int0_0_addr0 = i01_out;
        end else if((~(par_done_reg6_out | tmp_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            tmp_int0_0_addr0 = i00_out;
        end else tmp_int0_0_addr0 = 4'd0;
        if((((fsm7_out == 32'd5) & ~tmp_int0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            tmp_int0_0_addr1 = j01_out;
        end else if((~(par_done_reg6_out | tmp_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            tmp_int0_0_addr1 = j00_out;
        end else tmp_int0_0_addr1 = 4'd0;
        tmp_int0_0_clk = clk;
        if((((fsm7_out == 32'd5) & ~tmp_int0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            tmp_int0_0_write_data = tmp_sh_read0_0_out;
        end else tmp_int0_0_write_data = 32'd0;
        if((((fsm7_out == 32'd5) & ~tmp_int0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            tmp_int0_0_write_en = 1'd1;
        end else tmp_int0_0_write_en = 1'd0;
        if((((fsm_out == 32'd6) & ~j00_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            add0_left = j00_out;
        end else if((((fsm0_out == 32'd2) & ~i00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            add0_left = i00_out;
        end else if((((fsm1_out == 32'd5) & ~k0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            add0_left = k0_out;
        end else if((((fsm2_out == 32'd3) & ~j0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            add0_left = j0_out;
        end else if((((fsm3_out == 32'd2) & ~i0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            add0_left = i0_out;
        end else if((((fsm4_out == 32'd4) & ~k10_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            add0_left = k10_out;
        end else if((((fsm5_out == 32'd6) & ~j10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            add0_left = j10_out;
        end else if((((fsm6_out == 32'd2) & ~i10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            add0_left = i10_out;
        end else if((((fsm7_out == 32'd6) & ~j01_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            add0_left = j01_out;
        end else if((((fsm8_out == 32'd2) & ~i01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            add0_left = i01_out;
        end else add0_left = 4'd0;
        if((((fsm_out == 32'd6) & ~j00_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            add0_right = const14_out;
        end else if((((fsm0_out == 32'd2) & ~i00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            add0_right = const14_out;
        end else if((((fsm1_out == 32'd5) & ~k0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            add0_right = const14_out;
        end else if((((fsm2_out == 32'd3) & ~j0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            add0_right = const14_out;
        end else if((((fsm3_out == 32'd2) & ~i0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            add0_right = const14_out;
        end else if((((fsm4_out == 32'd4) & ~k10_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            add0_right = const14_out;
        end else if((((fsm5_out == 32'd6) & ~j10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            add0_right = const14_out;
        end else if((((fsm6_out == 32'd2) & ~i10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            add0_right = const14_out;
        end else if((((fsm7_out == 32'd6) & ~j01_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            add0_right = const14_out;
        end else if((((fsm8_out == 32'd2) & ~i01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            add0_right = const14_out;
        end else add0_right = 4'd0;
        if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            add2_left = tmp0_0_read_data;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            add2_left = D0_0_read_data;
        end else add2_left = 32'd0;
        if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            add2_right = v_0_out;
        end else if((((fsm4_out == 32'd3) & ~D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            add2_right = v1_0_out;
        end else add2_right = 32'd0;
        alpha_int_read0_0_clk = clk;
        if((~(par_done_reg7_out | alpha_int_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            alpha_int_read0_0_in = alpha_int0_read_data;
        end else alpha_int_read0_0_in = 32'd0;
        if((~(par_done_reg7_out | alpha_int_read0_0_done) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            alpha_int_read0_0_write_en = 1'd1;
        end else alpha_int_read0_0_write_en = 1'd0;
        beta_int_read0_0_clk = clk;
        if((((fsm5_out == 32'd1) & ~beta_int_read0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            beta_int_read0_0_in = beta_int0_read_data;
        end else beta_int_read0_0_in = 32'd0;
        if((((fsm5_out == 32'd1) & ~beta_int_read0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            beta_int_read0_0_write_en = 1'd1;
        end else beta_int_read0_0_write_en = 1'd0;
        bin_read0_0_clk = clk;
        if((((fsm1_out == 32'd1) & ~bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read0_0_in = mult_pipe0_out;
        end else bin_read0_0_in = 32'd0;
        if((((fsm1_out == 32'd1) & ~bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read0_0_write_en = mult_pipe0_done;
        end else bin_read0_0_write_en = 1'd0;
        bin_read1_0_clk = clk;
        if((((fsm1_out == 32'd2) & ~bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read1_0_in = mult_pipe1_out;
        end else bin_read1_0_in = 32'd0;
        if((((fsm1_out == 32'd2) & ~bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            bin_read1_0_write_en = mult_pipe1_done;
        end else bin_read1_0_write_en = 1'd0;
        bin_read2_0_clk = clk;
        if((((fsm5_out == 32'd2) & ~bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            bin_read2_0_in = mult_pipe2_out;
        end else bin_read2_0_in = 32'd0;
        if((((fsm5_out == 32'd2) & ~bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            bin_read2_0_write_en = mult_pipe2_done;
        end else bin_read2_0_write_en = 1'd0;
        bin_read3_0_clk = clk;
        if((((fsm4_out == 32'd1) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            bin_read3_0_in = mult_pipe3_out;
        end else bin_read3_0_in = 32'd0;
        if((((fsm4_out == 32'd1) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            bin_read3_0_write_en = mult_pipe3_done;
        end else bin_read3_0_write_en = 1'd0;
        cond_computed_clk = clk;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_computed_in = 1'd1;
        end else if((((cond_stored_out & cond_computed_out) & (fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_computed_in = 1'd0;
        end else if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_computed_in = 1'd0;
        end else cond_computed_in = 1'd0;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_computed_write_en = 1'd1;
        end else if((((cond_stored_out & cond_computed_out) & (fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_computed_write_en = 1'd1;
        end else if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_computed_write_en = 1'd1;
        end else cond_computed_write_en = 1'd0;
        cond_computed0_clk = clk;
        if((((~cond_computed0_out & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_computed0_in = 1'd1;
        end else if((((cond_stored0_out & cond_computed0_out) & (fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_computed0_in = 1'd0;
        end else if(((cond_computed0_out & ~cond_stored0_out) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_computed0_in = 1'd0;
        end else cond_computed0_in = 1'd0;
        if((((~cond_computed0_out & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_computed0_write_en = 1'd1;
        end else if((((cond_stored0_out & cond_computed0_out) & (fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_computed0_write_en = 1'd1;
        end else if(((cond_computed0_out & ~cond_stored0_out) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_computed0_write_en = 1'd1;
        end else cond_computed0_write_en = 1'd0;
        cond_computed1_clk = clk;
        if((((~cond_computed1_out & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_computed1_in = 1'd1;
        end else if((((cond_stored1_out & cond_computed1_out) & (fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_computed1_in = 1'd0;
        end else if(((cond_computed1_out & ~cond_stored1_out) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_computed1_in = 1'd0;
        end else cond_computed1_in = 1'd0;
        if((((~cond_computed1_out & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_computed1_write_en = 1'd1;
        end else if((((cond_stored1_out & cond_computed1_out) & (fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_computed1_write_en = 1'd1;
        end else if(((cond_computed1_out & ~cond_stored1_out) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_computed1_write_en = 1'd1;
        end else cond_computed1_write_en = 1'd0;
        cond_computed2_clk = clk;
        if((((~cond_computed2_out & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_in = 1'd1;
        end else if((((cond_stored2_out & cond_computed2_out) & (fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_in = 1'd0;
        end else if(((cond_computed2_out & ~cond_stored2_out) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_in = 1'd0;
        end else cond_computed2_in = 1'd0;
        if((((~cond_computed2_out & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_write_en = 1'd1;
        end else if((((cond_stored2_out & cond_computed2_out) & (fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_write_en = 1'd1;
        end else if(((cond_computed2_out & ~cond_stored2_out) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_computed2_write_en = 1'd1;
        end else cond_computed2_write_en = 1'd0;
        cond_computed3_clk = clk;
        if((((~cond_computed3_out & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_in = 1'd1;
        end else if((((cond_stored3_out & cond_computed3_out) & (fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_in = 1'd0;
        end else if(((cond_computed3_out & ~cond_stored3_out) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_in = 1'd0;
        end else cond_computed3_in = 1'd0;
        if((((~cond_computed3_out & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_write_en = 1'd1;
        end else if((((cond_stored3_out & cond_computed3_out) & (fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_write_en = 1'd1;
        end else if(((cond_computed3_out & ~cond_stored3_out) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_computed3_write_en = 1'd1;
        end else cond_computed3_write_en = 1'd0;
        cond_computed4_clk = clk;
        if((((~cond_computed4_out & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) & 1'b1) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_computed4_in = 1'd1;
        end else if((((cond_stored4_out & cond_computed4_out) & (fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_computed4_in = 1'd0;
        end else if(((cond_computed4_out & ~cond_stored4_out) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_computed4_in = 1'd0;
        end else cond_computed4_in = 1'd0;
        if((((~cond_computed4_out & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) & 1'b1) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_computed4_write_en = 1'd1;
        end else if((((cond_stored4_out & cond_computed4_out) & (fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_computed4_write_en = 1'd1;
        end else if(((cond_computed4_out & ~cond_stored4_out) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_computed4_write_en = 1'd1;
        end else cond_computed4_write_en = 1'd0;
        cond_computed5_clk = clk;
        if((((~cond_computed5_out & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_computed5_in = 1'd1;
        end else if((((cond_stored5_out & cond_computed5_out) & (fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_computed5_in = 1'd0;
        end else if(((cond_computed5_out & ~cond_stored5_out) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_computed5_in = 1'd0;
        end else cond_computed5_in = 1'd0;
        if((((~cond_computed5_out & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_computed5_write_en = 1'd1;
        end else if((((cond_stored5_out & cond_computed5_out) & (fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_computed5_write_en = 1'd1;
        end else if(((cond_computed5_out & ~cond_stored5_out) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_computed5_write_en = 1'd1;
        end else cond_computed5_write_en = 1'd0;
        cond_computed6_clk = clk;
        if((((~cond_computed6_out & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_in = 1'd1;
        end else if((((cond_stored6_out & cond_computed6_out) & (fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_in = 1'd0;
        end else if(((cond_computed6_out & ~cond_stored6_out) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_in = 1'd0;
        end else cond_computed6_in = 1'd0;
        if((((~cond_computed6_out & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_write_en = 1'd1;
        end else if((((cond_stored6_out & cond_computed6_out) & (fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_write_en = 1'd1;
        end else if(((cond_computed6_out & ~cond_stored6_out) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_computed6_write_en = 1'd1;
        end else cond_computed6_write_en = 1'd0;
        cond_computed7_clk = clk;
        if((((~cond_computed7_out & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_in = 1'd1;
        end else if((((cond_stored7_out & cond_computed7_out) & (fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_in = 1'd0;
        end else if(((cond_computed7_out & ~cond_stored7_out) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_in = 1'd0;
        end else cond_computed7_in = 1'd0;
        if((((~cond_computed7_out & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_write_en = 1'd1;
        end else if((((cond_stored7_out & cond_computed7_out) & (fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_write_en = 1'd1;
        end else if(((cond_computed7_out & ~cond_stored7_out) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_computed7_write_en = 1'd1;
        end else cond_computed7_write_en = 1'd0;
        cond_computed8_clk = clk;
        if((((~cond_computed8_out & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_in = 1'd1;
        end else if((((cond_stored8_out & cond_computed8_out) & (fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_in = 1'd0;
        end else if(((cond_computed8_out & ~cond_stored8_out) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_in = 1'd0;
        end else cond_computed8_in = 1'd0;
        if((((~cond_computed8_out & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_write_en = 1'd1;
        end else if((((cond_stored8_out & cond_computed8_out) & (fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_write_en = 1'd1;
        end else if(((cond_computed8_out & ~cond_stored8_out) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_computed8_write_en = 1'd1;
        end else cond_computed8_write_en = 1'd0;
        cond_stored_clk = clk;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_stored_in = le0_out;
        end else cond_stored_in = 1'd0;
        if((((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) & 1'b1) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            cond_stored_write_en = 1'd1;
        end else cond_stored_write_en = 1'd0;
        cond_stored0_clk = clk;
        if((((~cond_computed0_out & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_stored0_in = le0_out;
        end else cond_stored0_in = 1'd0;
        if((((~cond_computed0_out & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            cond_stored0_write_en = 1'd1;
        end else cond_stored0_write_en = 1'd0;
        cond_stored1_clk = clk;
        if((((~cond_computed1_out & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_stored1_in = le0_out;
        end else cond_stored1_in = 1'd0;
        if((((~cond_computed1_out & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) & 1'b1) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            cond_stored1_write_en = 1'd1;
        end else cond_stored1_write_en = 1'd0;
        cond_stored2_clk = clk;
        if((((~cond_computed2_out & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_stored2_in = le0_out;
        end else cond_stored2_in = 1'd0;
        if((((~cond_computed2_out & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) & 1'b1) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            cond_stored2_write_en = 1'd1;
        end else cond_stored2_write_en = 1'd0;
        cond_stored3_clk = clk;
        if((((~cond_computed3_out & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_stored3_in = le0_out;
        end else cond_stored3_in = 1'd0;
        if((((~cond_computed3_out & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            cond_stored3_write_en = 1'd1;
        end else cond_stored3_write_en = 1'd0;
        cond_stored4_clk = clk;
        if((((~cond_computed4_out & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) & 1'b1) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_stored4_in = le0_out;
        end else cond_stored4_in = 1'd0;
        if((((~cond_computed4_out & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) & 1'b1) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            cond_stored4_write_en = 1'd1;
        end else cond_stored4_write_en = 1'd0;
        cond_stored5_clk = clk;
        if((((~cond_computed5_out & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_stored5_in = le0_out;
        end else cond_stored5_in = 1'd0;
        if((((~cond_computed5_out & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) & 1'b1) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            cond_stored5_write_en = 1'd1;
        end else cond_stored5_write_en = 1'd0;
        cond_stored6_clk = clk;
        if((((~cond_computed6_out & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_stored6_in = le0_out;
        end else cond_stored6_in = 1'd0;
        if((((~cond_computed6_out & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            cond_stored6_write_en = 1'd1;
        end else cond_stored6_write_en = 1'd0;
        cond_stored7_clk = clk;
        if((((~cond_computed7_out & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_stored7_in = le0_out;
        end else cond_stored7_in = 1'd0;
        if((((~cond_computed7_out & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) & 1'b1) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            cond_stored7_write_en = 1'd1;
        end else cond_stored7_write_en = 1'd0;
        cond_stored8_clk = clk;
        if((((~cond_computed8_out & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_stored8_in = le0_out;
        end else cond_stored8_in = 1'd0;
        if((((~cond_computed8_out & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))) & 1'b1) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            cond_stored8_write_en = 1'd1;
        end else cond_stored8_write_en = 1'd0;
        d_tmp_0_clk = clk;
        if((((fsm5_out == 32'd0) & ~d_tmp_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            d_tmp_0_in = D0_0_read_data;
        end else d_tmp_0_in = 32'd0;
        if((((fsm5_out == 32'd0) & ~d_tmp_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            d_tmp_0_write_en = 1'd1;
        end else d_tmp_0_write_en = 1'd0;
        done_reg_clk = clk;
        if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            done_reg_in = 1'd1;
        end else if(done_reg_out) begin
            done_reg_in = 1'd0;
        end else done_reg_in = 1'd0;
        if(((cond_computed_out & ~cond_stored_out) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            done_reg_write_en = 1'd1;
        end else if(done_reg_out) begin
            done_reg_write_en = 1'd1;
        end else done_reg_write_en = 1'd0;
        done_reg0_clk = clk;
        if(((cond_computed0_out & ~cond_stored0_out) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            done_reg0_in = 1'd1;
        end else if(done_reg0_out) begin
            done_reg0_in = 1'd0;
        end else done_reg0_in = 1'd0;
        if(((cond_computed0_out & ~cond_stored0_out) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            done_reg0_write_en = 1'd1;
        end else if(done_reg0_out) begin
            done_reg0_write_en = 1'd1;
        end else done_reg0_write_en = 1'd0;
        done_reg1_clk = clk;
        if(((cond_computed1_out & ~cond_stored1_out) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            done_reg1_in = 1'd1;
        end else if(done_reg1_out) begin
            done_reg1_in = 1'd0;
        end else done_reg1_in = 1'd0;
        if(((cond_computed1_out & ~cond_stored1_out) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            done_reg1_write_en = 1'd1;
        end else if(done_reg1_out) begin
            done_reg1_write_en = 1'd1;
        end else done_reg1_write_en = 1'd0;
        done_reg2_clk = clk;
        if(((cond_computed2_out & ~cond_stored2_out) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            done_reg2_in = 1'd1;
        end else if(done_reg2_out) begin
            done_reg2_in = 1'd0;
        end else done_reg2_in = 1'd0;
        if(((cond_computed2_out & ~cond_stored2_out) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            done_reg2_write_en = 1'd1;
        end else if(done_reg2_out) begin
            done_reg2_write_en = 1'd1;
        end else done_reg2_write_en = 1'd0;
        done_reg3_clk = clk;
        if(((cond_computed3_out & ~cond_stored3_out) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            done_reg3_in = 1'd1;
        end else if(done_reg3_out) begin
            done_reg3_in = 1'd0;
        end else done_reg3_in = 1'd0;
        if(((cond_computed3_out & ~cond_stored3_out) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            done_reg3_write_en = 1'd1;
        end else if(done_reg3_out) begin
            done_reg3_write_en = 1'd1;
        end else done_reg3_write_en = 1'd0;
        done_reg4_clk = clk;
        if(((cond_computed4_out & ~cond_stored4_out) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            done_reg4_in = 1'd1;
        end else if(done_reg4_out) begin
            done_reg4_in = 1'd0;
        end else done_reg4_in = 1'd0;
        if(((cond_computed4_out & ~cond_stored4_out) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            done_reg4_write_en = 1'd1;
        end else if(done_reg4_out) begin
            done_reg4_write_en = 1'd1;
        end else done_reg4_write_en = 1'd0;
        done_reg5_clk = clk;
        if(((cond_computed5_out & ~cond_stored5_out) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            done_reg5_in = 1'd1;
        end else if(done_reg5_out) begin
            done_reg5_in = 1'd0;
        end else done_reg5_in = 1'd0;
        if(((cond_computed5_out & ~cond_stored5_out) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            done_reg5_write_en = 1'd1;
        end else if(done_reg5_out) begin
            done_reg5_write_en = 1'd1;
        end else done_reg5_write_en = 1'd0;
        done_reg6_clk = clk;
        if(((cond_computed6_out & ~cond_stored6_out) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            done_reg6_in = 1'd1;
        end else if(done_reg6_out) begin
            done_reg6_in = 1'd0;
        end else done_reg6_in = 1'd0;
        if(((cond_computed6_out & ~cond_stored6_out) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            done_reg6_write_en = 1'd1;
        end else if(done_reg6_out) begin
            done_reg6_write_en = 1'd1;
        end else done_reg6_write_en = 1'd0;
        done_reg7_clk = clk;
        if(((cond_computed7_out & ~cond_stored7_out) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            done_reg7_in = 1'd1;
        end else if(done_reg7_out) begin
            done_reg7_in = 1'd0;
        end else done_reg7_in = 1'd0;
        if(((cond_computed7_out & ~cond_stored7_out) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            done_reg7_write_en = 1'd1;
        end else if(done_reg7_out) begin
            done_reg7_write_en = 1'd1;
        end else done_reg7_write_en = 1'd0;
        done_reg8_clk = clk;
        if(((cond_computed8_out & ~cond_stored8_out) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            done_reg8_in = 1'd1;
        end else if(done_reg8_out) begin
            done_reg8_in = 1'd0;
        end else done_reg8_in = 1'd0;
        if(((cond_computed8_out & ~cond_stored8_out) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            done_reg8_write_en = 1'd1;
        end else if(done_reg8_out) begin
            done_reg8_write_en = 1'd1;
        end else done_reg8_write_en = 1'd0;
        fsm_clk = clk;
        if((((fsm_out == 32'd0) & A_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd1;
        end else if((((fsm_out == 32'd1) & par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd2;
        end else if((((fsm_out == 32'd2) & par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd3;
        end else if((((fsm_out == 32'd3) & par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd4;
        end else if((((fsm_out == 32'd4) & par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd5;
        end else if((((fsm_out == 32'd5) & tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd6;
        end else if((((fsm_out == 32'd6) & j00_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_in = 32'd7;
        end else if((fsm_out == 32'd7)) begin
            fsm_in = 32'd0;
        end else fsm_in = 32'd0;
        if((((fsm_out == 32'd0) & A_int_read0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd1) & par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd2) & par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd3) & par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd4) & par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd5) & tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((((fsm_out == 32'd6) & j00_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            fsm_write_en = 1'd1;
        end else if((fsm_out == 32'd7)) begin
            fsm_write_en = 1'd1;
        end else fsm_write_en = 1'd0;
        fsm0_clk = clk;
        if((((fsm0_out == 32'd0) & j00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            fsm0_in = 32'd1;
        end else if((((fsm0_out == 32'd1) & done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            fsm0_in = 32'd2;
        end else if((((fsm0_out == 32'd2) & i00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            fsm0_in = 32'd3;
        end else if((fsm0_out == 32'd3)) begin
            fsm0_in = 32'd0;
        end else fsm0_in = 32'd0;
        if((((fsm0_out == 32'd0) & j00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            fsm0_write_en = 1'd1;
        end else if((((fsm0_out == 32'd1) & done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            fsm0_write_en = 1'd1;
        end else if((((fsm0_out == 32'd2) & i00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            fsm0_write_en = 1'd1;
        end else if((fsm0_out == 32'd3)) begin
            fsm0_write_en = 1'd1;
        end else fsm0_write_en = 1'd0;
        fsm1_clk = clk;
        if((((fsm1_out == 32'd0) & par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_in = 32'd1;
        end else if((((fsm1_out == 32'd1) & bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_in = 32'd2;
        end else if((((fsm1_out == 32'd2) & bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_in = 32'd3;
        end else if((((fsm1_out == 32'd3) & v_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_in = 32'd4;
        end else if((((fsm1_out == 32'd4) & tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_in = 32'd5;
        end else if((((fsm1_out == 32'd5) & k0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_in = 32'd6;
        end else if((fsm1_out == 32'd6)) begin
            fsm1_in = 32'd0;
        end else fsm1_in = 32'd0;
        if((((fsm1_out == 32'd0) & par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd1) & bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd2) & bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd3) & v_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd4) & tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((((fsm1_out == 32'd5) & k0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            fsm1_write_en = 1'd1;
        end else if((fsm1_out == 32'd6)) begin
            fsm1_write_en = 1'd1;
        end else fsm1_write_en = 1'd0;
        fsm2_clk = clk;
        if((((fsm2_out == 32'd0) & tmp0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_in = 32'd1;
        end else if((((fsm2_out == 32'd1) & k0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_in = 32'd2;
        end else if((((fsm2_out == 32'd2) & done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_in = 32'd3;
        end else if((((fsm2_out == 32'd3) & j0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_in = 32'd4;
        end else if((fsm2_out == 32'd4)) begin
            fsm2_in = 32'd0;
        end else fsm2_in = 32'd0;
        if((((fsm2_out == 32'd0) & tmp0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((((fsm2_out == 32'd1) & k0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((((fsm2_out == 32'd2) & done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((((fsm2_out == 32'd3) & j0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            fsm2_write_en = 1'd1;
        end else if((fsm2_out == 32'd4)) begin
            fsm2_write_en = 1'd1;
        end else fsm2_write_en = 1'd0;
        fsm3_clk = clk;
        if((((fsm3_out == 32'd0) & j0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            fsm3_in = 32'd1;
        end else if((((fsm3_out == 32'd1) & done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            fsm3_in = 32'd2;
        end else if((((fsm3_out == 32'd2) & i0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            fsm3_in = 32'd3;
        end else if((fsm3_out == 32'd3)) begin
            fsm3_in = 32'd0;
        end else fsm3_in = 32'd0;
        if((((fsm3_out == 32'd0) & j0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            fsm3_write_en = 1'd1;
        end else if((((fsm3_out == 32'd1) & done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            fsm3_write_en = 1'd1;
        end else if((((fsm3_out == 32'd2) & i0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            fsm3_write_en = 1'd1;
        end else if((fsm3_out == 32'd3)) begin
            fsm3_write_en = 1'd1;
        end else fsm3_write_en = 1'd0;
        fsm4_clk = clk;
        if((((fsm4_out == 32'd0) & par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_in = 32'd1;
        end else if((((fsm4_out == 32'd1) & bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_in = 32'd2;
        end else if((((fsm4_out == 32'd2) & v1_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_in = 32'd3;
        end else if((((fsm4_out == 32'd3) & D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_in = 32'd4;
        end else if((((fsm4_out == 32'd4) & k10_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_in = 32'd5;
        end else if((fsm4_out == 32'd5)) begin
            fsm4_in = 32'd0;
        end else fsm4_in = 32'd0;
        if((((fsm4_out == 32'd0) & par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((((fsm4_out == 32'd1) & bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((((fsm4_out == 32'd2) & v1_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((((fsm4_out == 32'd3) & D0_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((((fsm4_out == 32'd4) & k10_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            fsm4_write_en = 1'd1;
        end else if((fsm4_out == 32'd5)) begin
            fsm4_write_en = 1'd1;
        end else fsm4_write_en = 1'd0;
        fsm5_clk = clk;
        if((((fsm5_out == 32'd0) & d_tmp_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd1;
        end else if((((fsm5_out == 32'd1) & beta_int_read0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd2;
        end else if((((fsm5_out == 32'd2) & bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd3;
        end else if((((fsm5_out == 32'd3) & D0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd4;
        end else if((((fsm5_out == 32'd4) & k10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd5;
        end else if((((fsm5_out == 32'd5) & done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd6;
        end else if((((fsm5_out == 32'd6) & j10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_in = 32'd7;
        end else if((fsm5_out == 32'd7)) begin
            fsm5_in = 32'd0;
        end else fsm5_in = 32'd0;
        if((((fsm5_out == 32'd0) & d_tmp_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd1) & beta_int_read0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd2) & bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd3) & D0_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd4) & k10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd5) & done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((((fsm5_out == 32'd6) & j10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            fsm5_write_en = 1'd1;
        end else if((fsm5_out == 32'd7)) begin
            fsm5_write_en = 1'd1;
        end else fsm5_write_en = 1'd0;
        fsm6_clk = clk;
        if((((fsm6_out == 32'd0) & j10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            fsm6_in = 32'd1;
        end else if((((fsm6_out == 32'd1) & done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            fsm6_in = 32'd2;
        end else if((((fsm6_out == 32'd2) & i10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            fsm6_in = 32'd3;
        end else if((fsm6_out == 32'd3)) begin
            fsm6_in = 32'd0;
        end else fsm6_in = 32'd0;
        if((((fsm6_out == 32'd0) & j10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            fsm6_write_en = 1'd1;
        end else if((((fsm6_out == 32'd1) & done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            fsm6_write_en = 1'd1;
        end else if((((fsm6_out == 32'd2) & i10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            fsm6_write_en = 1'd1;
        end else if((fsm6_out == 32'd3)) begin
            fsm6_write_en = 1'd1;
        end else fsm6_write_en = 1'd0;
        fsm7_clk = clk;
        if((((fsm7_out == 32'd0) & A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd1;
        end else if((((fsm7_out == 32'd1) & par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd2;
        end else if((((fsm7_out == 32'd2) & par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd3;
        end else if((((fsm7_out == 32'd3) & par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd4;
        end else if((((fsm7_out == 32'd4) & par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd5;
        end else if((((fsm7_out == 32'd5) & tmp_int0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd6;
        end else if((((fsm7_out == 32'd6) & j01_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_in = 32'd7;
        end else if((fsm7_out == 32'd7)) begin
            fsm7_in = 32'd0;
        end else fsm7_in = 32'd0;
        if((((fsm7_out == 32'd0) & A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd1) & par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd2) & par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd3) & par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd4) & par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd5) & tmp_int0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((((fsm7_out == 32'd6) & j01_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            fsm7_write_en = 1'd1;
        end else if((fsm7_out == 32'd7)) begin
            fsm7_write_en = 1'd1;
        end else fsm7_write_en = 1'd0;
        fsm8_clk = clk;
        if((((fsm8_out == 32'd0) & j01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            fsm8_in = 32'd1;
        end else if((((fsm8_out == 32'd1) & done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            fsm8_in = 32'd2;
        end else if((((fsm8_out == 32'd2) & i01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            fsm8_in = 32'd3;
        end else if((fsm8_out == 32'd3)) begin
            fsm8_in = 32'd0;
        end else fsm8_in = 32'd0;
        if((((fsm8_out == 32'd0) & j01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            fsm8_write_en = 1'd1;
        end else if((((fsm8_out == 32'd1) & done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            fsm8_write_en = 1'd1;
        end else if((((fsm8_out == 32'd2) & i01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            fsm8_write_en = 1'd1;
        end else if((fsm8_out == 32'd3)) begin
            fsm8_write_en = 1'd1;
        end else fsm8_write_en = 1'd0;
        fsm9_clk = clk;
        if((((fsm9_out == 32'd0) & i00_done) & (go | go))) begin
            fsm9_in = 32'd1;
        end else if((((fsm9_out == 32'd1) & done_reg0_out) & (go | go))) begin
            fsm9_in = 32'd2;
        end else if((((fsm9_out == 32'd2) & i0_done) & (go | go))) begin
            fsm9_in = 32'd3;
        end else if((((fsm9_out == 32'd3) & done_reg3_out) & (go | go))) begin
            fsm9_in = 32'd4;
        end else if((((fsm9_out == 32'd4) & i10_done) & (go | go))) begin
            fsm9_in = 32'd5;
        end else if((((fsm9_out == 32'd5) & done_reg6_out) & (go | go))) begin
            fsm9_in = 32'd6;
        end else if((((fsm9_out == 32'd6) & i01_done) & (go | go))) begin
            fsm9_in = 32'd7;
        end else if((((fsm9_out == 32'd7) & done_reg8_out) & (go | go))) begin
            fsm9_in = 32'd8;
        end else if((fsm9_out == 32'd8)) begin
            fsm9_in = 32'd0;
        end else fsm9_in = 32'd0;
        if((((fsm9_out == 32'd0) & i00_done) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd1) & done_reg0_out) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd2) & i0_done) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd3) & done_reg3_out) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd4) & i10_done) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd5) & done_reg6_out) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd6) & i01_done) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((((fsm9_out == 32'd7) & done_reg8_out) & (go | go))) begin
            fsm9_write_en = 1'd1;
        end else if((fsm9_out == 32'd8)) begin
            fsm9_write_en = 1'd1;
        end else fsm9_write_en = 1'd0;
        i0_clk = clk;
        if((((fsm9_out == 32'd2) & ~i0_done) & (go | go))) begin
            i0_in = const0_out;
        end else if((((fsm3_out == 32'd2) & ~i0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            i0_in = add0_out;
        end else i0_in = 4'd0;
        if((((fsm9_out == 32'd2) & ~i0_done) & (go | go))) begin
            i0_write_en = 1'd1;
        end else if((((fsm3_out == 32'd2) & ~i0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            i0_write_en = 1'd1;
        end else i0_write_en = 1'd0;
        i00_clk = clk;
        if((((fsm9_out == 32'd0) & ~i00_done) & (go | go))) begin
            i00_in = const0_out;
        end else if((((fsm0_out == 32'd2) & ~i00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            i00_in = add0_out;
        end else i00_in = 4'd0;
        if((((fsm9_out == 32'd0) & ~i00_done) & (go | go))) begin
            i00_write_en = 1'd1;
        end else if((((fsm0_out == 32'd2) & ~i00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            i00_write_en = 1'd1;
        end else i00_write_en = 1'd0;
        i01_clk = clk;
        if((((fsm9_out == 32'd6) & ~i01_done) & (go | go))) begin
            i01_in = const0_out;
        end else if((((fsm8_out == 32'd2) & ~i01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            i01_in = add0_out;
        end else i01_in = 4'd0;
        if((((fsm9_out == 32'd6) & ~i01_done) & (go | go))) begin
            i01_write_en = 1'd1;
        end else if((((fsm8_out == 32'd2) & ~i01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            i01_write_en = 1'd1;
        end else i01_write_en = 1'd0;
        i10_clk = clk;
        if((((fsm9_out == 32'd4) & ~i10_done) & (go | go))) begin
            i10_in = const0_out;
        end else if((((fsm6_out == 32'd2) & ~i10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            i10_in = add0_out;
        end else i10_in = 4'd0;
        if((((fsm9_out == 32'd4) & ~i10_done) & (go | go))) begin
            i10_write_en = 1'd1;
        end else if((((fsm6_out == 32'd2) & ~i10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            i10_write_en = 1'd1;
        end else i10_write_en = 1'd0;
        j0_clk = clk;
        if((((fsm3_out == 32'd0) & ~j0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            j0_in = const0_out;
        end else if((((fsm2_out == 32'd3) & ~j0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            j0_in = add0_out;
        end else j0_in = 4'd0;
        if((((fsm3_out == 32'd0) & ~j0_done) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))) begin
            j0_write_en = 1'd1;
        end else if((((fsm2_out == 32'd3) & ~j0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            j0_write_en = 1'd1;
        end else j0_write_en = 1'd0;
        j00_clk = clk;
        if((((fsm0_out == 32'd0) & ~j00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            j00_in = const0_out;
        end else if((((fsm_out == 32'd6) & ~j00_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            j00_in = add0_out;
        end else j00_in = 4'd0;
        if((((fsm0_out == 32'd0) & ~j00_done) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))) begin
            j00_write_en = 1'd1;
        end else if((((fsm_out == 32'd6) & ~j00_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            j00_write_en = 1'd1;
        end else j00_write_en = 1'd0;
        j01_clk = clk;
        if((((fsm8_out == 32'd0) & ~j01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            j01_in = const0_out;
        end else if((((fsm7_out == 32'd6) & ~j01_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            j01_in = add0_out;
        end else j01_in = 4'd0;
        if((((fsm8_out == 32'd0) & ~j01_done) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))) begin
            j01_write_en = 1'd1;
        end else if((((fsm7_out == 32'd6) & ~j01_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            j01_write_en = 1'd1;
        end else j01_write_en = 1'd0;
        j10_clk = clk;
        if((((fsm6_out == 32'd0) & ~j10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            j10_in = const0_out;
        end else if((((fsm5_out == 32'd6) & ~j10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            j10_in = add0_out;
        end else j10_in = 4'd0;
        if((((fsm6_out == 32'd0) & ~j10_done) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))) begin
            j10_write_en = 1'd1;
        end else if((((fsm5_out == 32'd6) & ~j10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            j10_write_en = 1'd1;
        end else j10_write_en = 1'd0;
        k0_clk = clk;
        if((((fsm2_out == 32'd1) & ~k0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            k0_in = const0_out;
        end else if((((fsm1_out == 32'd5) & ~k0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            k0_in = add0_out;
        end else k0_in = 4'd0;
        if((((fsm2_out == 32'd1) & ~k0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            k0_write_en = 1'd1;
        end else if((((fsm1_out == 32'd5) & ~k0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            k0_write_en = 1'd1;
        end else k0_write_en = 1'd0;
        k10_clk = clk;
        if((((fsm5_out == 32'd4) & ~k10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            k10_in = const0_out;
        end else if((((fsm4_out == 32'd4) & ~k10_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            k10_in = add0_out;
        end else k10_in = 4'd0;
        if((((fsm5_out == 32'd4) & ~k10_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            k10_write_en = 1'd1;
        end else if((((fsm4_out == 32'd4) & ~k10_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            k10_write_en = 1'd1;
        end else k10_write_en = 1'd0;
        if((~cond_computed0_out & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            le0_left = i00_out;
        end else if((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            le0_left = j00_out;
        end else if((~cond_computed3_out & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            le0_left = i0_out;
        end else if((~cond_computed2_out & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            le0_left = j0_out;
        end else if((~cond_computed1_out & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            le0_left = k0_out;
        end else if((~cond_computed6_out & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            le0_left = i10_out;
        end else if((~cond_computed5_out & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            le0_left = j10_out;
        end else if((~cond_computed4_out & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            le0_left = k10_out;
        end else if((~cond_computed8_out & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            le0_left = i01_out;
        end else if((~cond_computed7_out & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            le0_left = j01_out;
        end else le0_left = 4'd0;
        if((~cond_computed0_out & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))) begin
            le0_right = const1_out;
        end else if((~cond_computed_out & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))) begin
            le0_right = const1_out;
        end else if((~cond_computed3_out & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))) begin
            le0_right = const1_out;
        end else if((~cond_computed2_out & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))) begin
            le0_right = const1_out;
        end else if((~cond_computed1_out & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))) begin
            le0_right = const1_out;
        end else if((~cond_computed6_out & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))) begin
            le0_right = const1_out;
        end else if((~cond_computed5_out & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))) begin
            le0_right = const1_out;
        end else if((~cond_computed4_out & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            le0_right = const1_out;
        end else if((~cond_computed8_out & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))) begin
            le0_right = const1_out;
        end else if((~cond_computed7_out & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))) begin
            le0_right = const1_out;
        end else le0_right = 4'd0;
        mult_pipe0_clk = clk;
        if((~mult_pipe0_done & (((fsm1_out == 32'd1) & ~bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            mult_pipe0_go = 1'd1;
        end else mult_pipe0_go = 1'd0;
        if((((fsm1_out == 32'd1) & ~bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe0_left = alpha_int_read0_0_out;
        end else mult_pipe0_left = 32'd0;
        if((((fsm1_out == 32'd1) & ~bin_read0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe0_right = A_read0_0_out;
        end else mult_pipe0_right = 32'd0;
        mult_pipe1_clk = clk;
        if((~mult_pipe1_done & (((fsm1_out == 32'd2) & ~bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            mult_pipe1_go = 1'd1;
        end else mult_pipe1_go = 1'd0;
        if((((fsm1_out == 32'd2) & ~bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe1_left = bin_read0_0_out;
        end else mult_pipe1_left = 32'd0;
        if((((fsm1_out == 32'd2) & ~bin_read1_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            mult_pipe1_right = B_read0_0_out;
        end else mult_pipe1_right = 32'd0;
        mult_pipe2_clk = clk;
        if((~mult_pipe2_done & (((fsm5_out == 32'd2) & ~bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))) begin
            mult_pipe2_go = 1'd1;
        end else mult_pipe2_go = 1'd0;
        if((((fsm5_out == 32'd2) & ~bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            mult_pipe2_left = beta_int_read0_0_out;
        end else mult_pipe2_left = 32'd0;
        if((((fsm5_out == 32'd2) & ~bin_read2_0_done) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))) begin
            mult_pipe2_right = d_tmp_0_out;
        end else mult_pipe2_right = 32'd0;
        mult_pipe3_clk = clk;
        if((~mult_pipe3_done & (((fsm4_out == 32'd1) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            mult_pipe3_go = 1'd1;
        end else mult_pipe3_go = 1'd0;
        if((((fsm4_out == 32'd1) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            mult_pipe3_left = tmp_read0_0_out;
        end else mult_pipe3_left = 32'd0;
        if((((fsm4_out == 32'd1) & ~bin_read3_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            mult_pipe3_right = C_read0_0_out;
        end else mult_pipe3_right = 32'd0;
        par_done_reg_clk = clk;
        if((A0_0_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg_in = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg_in = 1'd0;
        end else par_done_reg_in = 1'd0;
        if((A0_0_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg_write_en = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg_write_en = 1'd1;
        end else par_done_reg_write_en = 1'd0;
        par_done_reg0_clk = clk;
        if((B_int_read0_0_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg0_in = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg0_in = 1'd0;
        end else par_done_reg0_in = 1'd0;
        if((B_int_read0_0_done & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg0_write_en = 1'd1;
        end else if(par_reset_out) begin
            par_done_reg0_write_en = 1'd1;
        end else par_done_reg0_write_en = 1'd0;
        par_done_reg1_clk = clk;
        if((B0_0_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg1_in = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg1_in = 1'd0;
        end else par_done_reg1_in = 1'd0;
        if((B0_0_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg1_write_en = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg1_write_en = 1'd1;
        end else par_done_reg1_write_en = 1'd0;
        par_done_reg10_clk = clk;
        if((tmp_read0_0_done & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            par_done_reg10_in = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg10_in = 1'd0;
        end else par_done_reg10_in = 1'd0;
        if((tmp_read0_0_done & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            par_done_reg10_write_en = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg10_write_en = 1'd1;
        end else par_done_reg10_write_en = 1'd0;
        par_done_reg11_clk = clk;
        if((C_read0_0_done & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            par_done_reg11_in = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg11_in = 1'd0;
        end else par_done_reg11_in = 1'd0;
        if((C_read0_0_done & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            par_done_reg11_write_en = 1'd1;
        end else if(par_reset4_out) begin
            par_done_reg11_write_en = 1'd1;
        end else par_done_reg11_write_en = 1'd0;
        par_done_reg12_clk = clk;
        if((A_int0_0_done & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg12_in = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg12_in = 1'd0;
        end else par_done_reg12_in = 1'd0;
        if((A_int0_0_done & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg12_write_en = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg12_write_en = 1'd1;
        end else par_done_reg12_write_en = 1'd0;
        par_done_reg13_clk = clk;
        if((B_sh_read0_0_done & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg13_in = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg13_in = 1'd0;
        end else par_done_reg13_in = 1'd0;
        if((B_sh_read0_0_done & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg13_write_en = 1'd1;
        end else if(par_reset5_out) begin
            par_done_reg13_write_en = 1'd1;
        end else par_done_reg13_write_en = 1'd0;
        par_done_reg14_clk = clk;
        if((B_int0_0_done & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg14_in = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg14_in = 1'd0;
        end else par_done_reg14_in = 1'd0;
        if((B_int0_0_done & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg14_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg14_write_en = 1'd1;
        end else par_done_reg14_write_en = 1'd0;
        par_done_reg15_clk = clk;
        if((C_sh_read0_0_done & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg15_in = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg15_in = 1'd0;
        end else par_done_reg15_in = 1'd0;
        if((C_sh_read0_0_done & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg15_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_done_reg15_write_en = 1'd1;
        end else par_done_reg15_write_en = 1'd0;
        par_done_reg16_clk = clk;
        if((C_int0_0_done & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg16_in = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg16_in = 1'd0;
        end else par_done_reg16_in = 1'd0;
        if((C_int0_0_done & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg16_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg16_write_en = 1'd1;
        end else par_done_reg16_write_en = 1'd0;
        par_done_reg17_clk = clk;
        if((D_sh_read0_0_done & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg17_in = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg17_in = 1'd0;
        end else par_done_reg17_in = 1'd0;
        if((D_sh_read0_0_done & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg17_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_done_reg17_write_en = 1'd1;
        end else par_done_reg17_write_en = 1'd0;
        par_done_reg18_clk = clk;
        if((D_int0_0_done & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg18_in = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg18_in = 1'd0;
        end else par_done_reg18_in = 1'd0;
        if((D_int0_0_done & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg18_write_en = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg18_write_en = 1'd1;
        end else par_done_reg18_write_en = 1'd0;
        par_done_reg19_clk = clk;
        if((tmp_sh_read0_0_done & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg19_in = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg19_in = 1'd0;
        end else par_done_reg19_in = 1'd0;
        if((tmp_sh_read0_0_done & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_done_reg19_write_en = 1'd1;
        end else if(par_reset8_out) begin
            par_done_reg19_write_en = 1'd1;
        end else par_done_reg19_write_en = 1'd0;
        par_done_reg2_clk = clk;
        if((C_int_read0_0_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg2_in = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg2_in = 1'd0;
        end else par_done_reg2_in = 1'd0;
        if((C_int_read0_0_done & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg2_write_en = 1'd1;
        end else if(par_reset0_out) begin
            par_done_reg2_write_en = 1'd1;
        end else par_done_reg2_write_en = 1'd0;
        par_done_reg3_clk = clk;
        if((C0_0_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg3_in = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg3_in = 1'd0;
        end else par_done_reg3_in = 1'd0;
        if((C0_0_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg3_write_en = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg3_write_en = 1'd1;
        end else par_done_reg3_write_en = 1'd0;
        par_done_reg4_clk = clk;
        if((D_int_read0_0_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg4_in = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg4_in = 1'd0;
        end else par_done_reg4_in = 1'd0;
        if((D_int_read0_0_done & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg4_write_en = 1'd1;
        end else if(par_reset1_out) begin
            par_done_reg4_write_en = 1'd1;
        end else par_done_reg4_write_en = 1'd0;
        par_done_reg5_clk = clk;
        if((D0_0_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg5_in = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg5_in = 1'd0;
        end else par_done_reg5_in = 1'd0;
        if((D0_0_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg5_write_en = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg5_write_en = 1'd1;
        end else par_done_reg5_write_en = 1'd0;
        par_done_reg6_clk = clk;
        if((tmp_int_read0_0_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg6_in = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg6_in = 1'd0;
        end else par_done_reg6_in = 1'd0;
        if((tmp_int_read0_0_done & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_done_reg6_write_en = 1'd1;
        end else if(par_reset2_out) begin
            par_done_reg6_write_en = 1'd1;
        end else par_done_reg6_write_en = 1'd0;
        par_done_reg7_clk = clk;
        if((alpha_int_read0_0_done & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_done_reg7_in = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg7_in = 1'd0;
        end else par_done_reg7_in = 1'd0;
        if((alpha_int_read0_0_done & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_done_reg7_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg7_write_en = 1'd1;
        end else par_done_reg7_write_en = 1'd0;
        par_done_reg8_clk = clk;
        if((A_read0_0_done & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_done_reg8_in = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg8_in = 1'd0;
        end else par_done_reg8_in = 1'd0;
        if((A_read0_0_done & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_done_reg8_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg8_write_en = 1'd1;
        end else par_done_reg8_write_en = 1'd0;
        par_done_reg9_clk = clk;
        if((B_read0_0_done & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_done_reg9_in = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg9_in = 1'd0;
        end else par_done_reg9_in = 1'd0;
        if((B_read0_0_done & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_done_reg9_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_done_reg9_write_en = 1'd1;
        end else par_done_reg9_write_en = 1'd0;
        par_reset_clk = clk;
        if(((par_done_reg_out & par_done_reg0_out) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset_in = 1'd1;
        end else if(par_reset_out) begin
            par_reset_in = 1'd0;
        end else par_reset_in = 1'd0;
        if(((par_done_reg_out & par_done_reg0_out) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset_write_en = 1'd1;
        end else if(par_reset_out) begin
            par_reset_write_en = 1'd1;
        end else par_reset_write_en = 1'd0;
        par_reset0_clk = clk;
        if(((par_done_reg1_out & par_done_reg2_out) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset0_in = 1'd1;
        end else if(par_reset0_out) begin
            par_reset0_in = 1'd0;
        end else par_reset0_in = 1'd0;
        if(((par_done_reg1_out & par_done_reg2_out) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset0_write_en = 1'd1;
        end else if(par_reset0_out) begin
            par_reset0_write_en = 1'd1;
        end else par_reset0_write_en = 1'd0;
        par_reset1_clk = clk;
        if(((par_done_reg3_out & par_done_reg4_out) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset1_in = 1'd1;
        end else if(par_reset1_out) begin
            par_reset1_in = 1'd0;
        end else par_reset1_in = 1'd0;
        if(((par_done_reg3_out & par_done_reg4_out) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset1_write_en = 1'd1;
        end else if(par_reset1_out) begin
            par_reset1_write_en = 1'd1;
        end else par_reset1_write_en = 1'd0;
        par_reset2_clk = clk;
        if(((par_done_reg5_out & par_done_reg6_out) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset2_in = 1'd1;
        end else if(par_reset2_out) begin
            par_reset2_in = 1'd0;
        end else par_reset2_in = 1'd0;
        if(((par_done_reg5_out & par_done_reg6_out) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            par_reset2_write_en = 1'd1;
        end else if(par_reset2_out) begin
            par_reset2_write_en = 1'd1;
        end else par_reset2_write_en = 1'd0;
        par_reset3_clk = clk;
        if((((par_done_reg7_out & par_done_reg8_out) & par_done_reg9_out) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_reset3_in = 1'd1;
        end else if(par_reset3_out) begin
            par_reset3_in = 1'd0;
        end else par_reset3_in = 1'd0;
        if((((par_done_reg7_out & par_done_reg8_out) & par_done_reg9_out) & (((fsm1_out == 32'd0) & ~par_reset3_out) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go)))))))))) begin
            par_reset3_write_en = 1'd1;
        end else if(par_reset3_out) begin
            par_reset3_write_en = 1'd1;
        end else par_reset3_write_en = 1'd0;
        par_reset4_clk = clk;
        if(((par_done_reg10_out & par_done_reg11_out) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            par_reset4_in = 1'd1;
        end else if(par_reset4_out) begin
            par_reset4_in = 1'd0;
        end else par_reset4_in = 1'd0;
        if(((par_done_reg10_out & par_done_reg11_out) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            par_reset4_write_en = 1'd1;
        end else if(par_reset4_out) begin
            par_reset4_write_en = 1'd1;
        end else par_reset4_write_en = 1'd0;
        par_reset5_clk = clk;
        if(((par_done_reg12_out & par_done_reg13_out) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset5_in = 1'd1;
        end else if(par_reset5_out) begin
            par_reset5_in = 1'd0;
        end else par_reset5_in = 1'd0;
        if(((par_done_reg12_out & par_done_reg13_out) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset5_write_en = 1'd1;
        end else if(par_reset5_out) begin
            par_reset5_write_en = 1'd1;
        end else par_reset5_write_en = 1'd0;
        par_reset6_clk = clk;
        if(((par_done_reg14_out & par_done_reg15_out) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset6_in = 1'd1;
        end else if(par_reset6_out) begin
            par_reset6_in = 1'd0;
        end else par_reset6_in = 1'd0;
        if(((par_done_reg14_out & par_done_reg15_out) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset6_write_en = 1'd1;
        end else if(par_reset6_out) begin
            par_reset6_write_en = 1'd1;
        end else par_reset6_write_en = 1'd0;
        par_reset7_clk = clk;
        if(((par_done_reg16_out & par_done_reg17_out) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset7_in = 1'd1;
        end else if(par_reset7_out) begin
            par_reset7_in = 1'd0;
        end else par_reset7_in = 1'd0;
        if(((par_done_reg16_out & par_done_reg17_out) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset7_write_en = 1'd1;
        end else if(par_reset7_out) begin
            par_reset7_write_en = 1'd1;
        end else par_reset7_write_en = 1'd0;
        par_reset8_clk = clk;
        if(((par_done_reg18_out & par_done_reg19_out) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset8_in = 1'd1;
        end else if(par_reset8_out) begin
            par_reset8_in = 1'd0;
        end else par_reset8_in = 1'd0;
        if(((par_done_reg18_out & par_done_reg19_out) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            par_reset8_write_en = 1'd1;
        end else if(par_reset8_out) begin
            par_reset8_write_en = 1'd1;
        end else par_reset8_write_en = 1'd0;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_left = j00_out;
        end else if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            rsh0_left = j01_out;
        end else if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_left = j00_out;
        end else if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_left = j01_out;
        end else if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_left = j01_out;
        end else if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_left = j01_out;
        end else if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_left = j01_out;
        end else if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_left = j00_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_left = j00_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            rsh0_left = j00_out;
        end else rsh0_left = 4'd0;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh0_right = const0_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            rsh0_right = const0_out;
        end else rsh0_right = 4'd0;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_left = i00_out;
        end else if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            rsh1_left = i01_out;
        end else if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_left = i00_out;
        end else if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_left = i01_out;
        end else if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_left = i01_out;
        end else if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_left = i01_out;
        end else if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_left = i01_out;
        end else if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_left = i00_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_left = i00_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            rsh1_left = i00_out;
        end else rsh1_left = 4'd0;
        if((~(par_done_reg_out | A0_0_done) & (((fsm_out == 32'd1) & ~par_reset_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((((fsm7_out == 32'd0) & ~A_sh_read0_0_done) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg1_out | B0_0_done) & (((fsm_out == 32'd2) & ~par_reset0_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg13_out | B_sh_read0_0_done) & (((fsm7_out == 32'd1) & ~par_reset5_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg15_out | C_sh_read0_0_done) & (((fsm7_out == 32'd2) & ~par_reset6_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg17_out | D_sh_read0_0_done) & (((fsm7_out == 32'd3) & ~par_reset7_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg3_out | C0_0_done) & (((fsm_out == 32'd3) & ~par_reset1_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((~(par_done_reg5_out | D0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            rsh1_right = const10_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            rsh1_right = const10_out;
        end else rsh1_right = 4'd0;
        if((((fsm2_out == 32'd0) & ~tmp0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            tmp0_0_addr0 = i0_out;
        end else if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            tmp0_0_addr0 = i0_out;
        end else if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            tmp0_0_addr0 = i0_out;
        end else if((~(par_done_reg10_out | tmp_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            tmp0_0_addr0 = i10_out;
        end else if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            tmp0_0_addr0 = rsh1_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            tmp0_0_addr0 = rsh1_out;
        end else tmp0_0_addr0 = 4'd0;
        if((((fsm2_out == 32'd0) & ~tmp0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            tmp0_0_addr1 = j0_out;
        end else if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            tmp0_0_addr1 = j0_out;
        end else if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            tmp0_0_addr1 = j0_out;
        end else if((~(par_done_reg10_out | tmp_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            tmp0_0_addr1 = k10_out;
        end else if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            tmp0_0_addr1 = rsh0_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            tmp0_0_addr1 = rsh0_out;
        end else tmp0_0_addr1 = 4'd0;
        tmp0_0_clk = clk;
        if((((fsm2_out == 32'd0) & ~tmp0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            tmp0_0_write_data = const20_out;
        end else if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            tmp0_0_write_data = add2_out;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            tmp0_0_write_data = tmp_int_read0_0_out;
        end else tmp0_0_write_data = 32'd0;
        if((((fsm2_out == 32'd0) & ~tmp0_0_done) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))) begin
            tmp0_0_write_en = 1'd1;
        end else if((((fsm1_out == 32'd4) & ~tmp0_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            tmp0_0_write_en = 1'd1;
        end else if((((fsm_out == 32'd5) & ~tmp0_0_done) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go))))))) begin
            tmp0_0_write_en = 1'd1;
        end else tmp0_0_write_en = 1'd0;
        tmp_int_read0_0_clk = clk;
        if((~(par_done_reg6_out | tmp_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            tmp_int_read0_0_in = tmp_int0_0_read_data;
        end else tmp_int_read0_0_in = 32'd0;
        if((~(par_done_reg6_out | tmp_int_read0_0_done) & (((fsm_out == 32'd4) & ~par_reset2_out) & (((cond_stored_out & cond_computed_out) & ~(fsm_out == 32'd7)) & (((fsm0_out == 32'd1) & ~done_reg_out) & (((cond_stored0_out & cond_computed0_out) & ~(fsm0_out == 32'd3)) & (((fsm9_out == 32'd1) & ~done_reg0_out) & (go | go)))))))) begin
            tmp_int_read0_0_write_en = 1'd1;
        end else tmp_int_read0_0_write_en = 1'd0;
        tmp_read0_0_clk = clk;
        if((~(par_done_reg10_out | tmp_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            tmp_read0_0_in = tmp0_0_read_data;
        end else tmp_read0_0_in = 32'd0;
        if((~(par_done_reg10_out | tmp_read0_0_done) & (((fsm4_out == 32'd0) & ~par_reset4_out) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go)))))))))) begin
            tmp_read0_0_write_en = 1'd1;
        end else tmp_read0_0_write_en = 1'd0;
        tmp_sh_read0_0_clk = clk;
        if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            tmp_sh_read0_0_in = tmp0_0_read_data;
        end else tmp_sh_read0_0_in = 32'd0;
        if((~(par_done_reg19_out | tmp_sh_read0_0_done) & (((fsm7_out == 32'd4) & ~par_reset8_out) & (((cond_stored7_out & cond_computed7_out) & ~(fsm7_out == 32'd7)) & (((fsm8_out == 32'd1) & ~done_reg7_out) & (((cond_stored8_out & cond_computed8_out) & ~(fsm8_out == 32'd3)) & (((fsm9_out == 32'd7) & ~done_reg8_out) & (go | go)))))))) begin
            tmp_sh_read0_0_write_en = 1'd1;
        end else tmp_sh_read0_0_write_en = 1'd0;
        v1_0_clk = clk;
        if((((fsm4_out == 32'd2) & ~v1_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            v1_0_in = bin_read3_0_out;
        end else v1_0_in = 32'd0;
        if((((fsm4_out == 32'd2) & ~v1_0_done) & (((cond_stored4_out & cond_computed4_out) & ~(fsm4_out == 32'd5)) & (((fsm5_out == 32'd5) & ~done_reg4_out) & (((cond_stored5_out & cond_computed5_out) & ~(fsm5_out == 32'd7)) & (((fsm6_out == 32'd1) & ~done_reg5_out) & (((cond_stored6_out & cond_computed6_out) & ~(fsm6_out == 32'd3)) & (((fsm9_out == 32'd5) & ~done_reg6_out) & (go | go))))))))) begin
            v1_0_write_en = 1'd1;
        end else v1_0_write_en = 1'd0;
        v_0_clk = clk;
        if((((fsm1_out == 32'd3) & ~v_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            v_0_in = bin_read1_0_out;
        end else v_0_in = 32'd0;
        if((((fsm1_out == 32'd3) & ~v_0_done) & (((cond_stored1_out & cond_computed1_out) & ~(fsm1_out == 32'd6)) & (((fsm2_out == 32'd2) & ~done_reg1_out) & (((cond_stored2_out & cond_computed2_out) & ~(fsm2_out == 32'd4)) & (((fsm3_out == 32'd1) & ~done_reg2_out) & (((cond_stored3_out & cond_computed3_out) & ~(fsm3_out == 32'd3)) & (((fsm9_out == 32'd3) & ~done_reg3_out) & (go | go))))))))) begin
            v_0_write_en = 1'd1;
        end else v_0_write_en = 1'd0;
    end
endmodule
